PK   �|�X�?p�Y  j�     cirkitFile.json�]m��6�+��`��H�6mq�M� ��ł����^˕�\��~���ږd�3LRnd���pH>�)�CԘ7vy�׍�{c�uU/�k"fѽi��f�i2�V���~o��>���?�������aU/�K
%%3"Ns�bnJ�T�X$9�ɥ��]]���}2;��S;ñs����8v�cW8v��vwc�J���Kbd�e�Ɔ�y�%L����X�`���NT]�D�B��<�9*64���Ds�����L�l��D����6�6ձQ�Ĳɬ�Xd�|��<-�D%6�DјSV�Y�t�uj|�SZd�b�j��2/�����Ն�ؤY+�2^���B �N10#8�IT�U�BՍ�s�i�H�B�.��(ҩQ�W�H�F�~�"Ez6��C�!�ǰ1�?��C�M������hŠ�"���@=Y �D�S�0�iH@4�a��F�C��qC5���*Tw��yڨ�B�T�Q��7f���� ��8/pJ#�<�?@����>�=@����>��اC�,��2�iR�L.ˡ�-LݸY���FN��/�D��
ӊ	�&Ȱ\
f���@��2_�T
��"���K[���n�i�蛤��� ��� Rh),�D�"%"E���H�aP�[��9FL_�$�Ĉ��m�(�����L���q�MYZ�L�p�׋�L��aX�$a#fbQ2��4�i ��0V��1�4��a1c�iSLà��A1�b(��b�,�Y��(�fy�E'E�g)䜳�&PO�Є��A����	h��t��9��#M�B��.4�_�Nkh�-�����u �c���B�.xɹ��\;���d��ip�+D߄A09y�3�9`^��"�b:�4]�[�=e~֭i-6󳴛�1d�/��H�A�� R� Rd)*�u���$|I��0 &aL�@���0	b�4�i �4�i�0(�aPLà��A1�b�,�Y�P"�Y�0(faP�΢���K9�p��p�/�l�����R�����-g~�R��kp�/��g~�R��ip�/�_�g~�	���kx�'��0 >�F�g~N�%h�/��p�3?x)��|��?ߵ�����x]�Y��j��n�0�-��]����_�6c|��u�3n��'t��P�0AU�p�U�ľ��<�IQ�	F�=�C	>v��A�5���?�
~��&z���D��/Y`^����noZc�7Σ�e1��^;�������4@:�  �] �n/�X�@���P�Oj�%<�gS � O*�%��i|w�����yz�i�bS-w�v�벌vG6U�=8p�<2��H~���H~��O��ɯ���4 =���+t(�B
�C�����Pos�����|F�H�DT?,p$o"ڄ�8��zS;(vP��a���k�)�S�!�XKL���b�ȰHdX$2t8�E"�"�a�ȰHd'���?���k�>�a�����aު�7��$��6|`���Hs0y���
�;'�>� ����o�c�O8 �V?
]hx��>�;Ack�����$���"�`!KN9+�>?l
�7����{�j>p$��� Ob���t���O�@ܽ�~�{�L�V���c���c���m�Ӊt����6�v.�̓.�%��$v�L'��z����sP�A=��sP�A=��s�N��<��s��^!��?l�c�8��A���	A�S���=��M��m=V�����5u/Η9=2����pJ�A(�vG���!��#�;v2���;ː'Q�Nw��p��g�n6C�W�$����+Ʒb��w�c��	���bz� �?��0�]tA���D�����64�]�m�m�m�m��ۢtX$�ErX��E�`f���7W��4�xJY�-�u����]��0�q�>t�^6��6me�(�a����0�:�mS-w�,̓��Kg����O�um�]�YV�������߾X>sr���,���m�[�����=k쟛��Et�6��`������)���4�7h�_s��U�}I�k.�\̘dsI%q ���M��s�y�#��Te��#D��P��٤���3J�^����b�Y�B��,�^(��EuS9)��0j���[/�j���kN�k�I*�8�q)��v��39Y4¥�$�cѐK$�u��aq%��s�����D�q>.'��=�������:NF�qufL����I:���jg���k��9	�	T��@�9	�?֏���}4��3�W.����c��>�,J���z�<�u�^	��I�x�{�/�Ӿh؛��.�����zQ�f�ᦳ�7��M��ö��M4����{b(e):NJ����]DUg&s�ψNs���w�E��?ڇ�󞗔��"W1)I�ySg�X'$�sg㤲E���������,.2��X@�`��c�]HER�2����/W�v���2-	wj�4w���\��Gr�'R��r�7p�|���"~v}r�h˟Z��Z����R*nbZ�XÅ7.̐��%�D��jj�AW<3MS�/Vv�'Er-h��XQ^ļp!jf]�&�M��:�Ɉ�g�zm��q� 3AT�l�Z�]wi���s�RUd9��v��ne�����=�g�s5�{�ӟٲ���y�\?TySw����<�d��eݴ�Ec��m��Ygge��#�;�}�eJ4/�XȔ������c��4sNP1]NAL�܅�$��"�ݹ�6&���HR�l��1�1�I]�I�9>M�X'n,I�Tʉ�ѩ����׹.cA��zFb]
g�b�8/K�8���x����jm���o��ps������+W���z��%W����6vv��W�fyU;w�ݿ���NТ���<�j9"��+kZ[,���5e6o;�tZ�%�������� ���;3G洋vn��⏪}�n���.����bH��_!x,L�l������xאЁ��
{k��(=�\��p�����٦nIE���M�MA
�;�v����$(e	'I�:O.�w�?$���]St2^�&�o#��?�>'��L�T�E`R�1f\#��5St;I��>}~��������X��_�n?~��k�
�]�q�y<,lnR)�w��J�{Ҳ�)+c�� ��v5��q����?Z�y�%%�'�͝�I���)�Z&��S�1%jN�[�?bo���s�4�z�M�&-努ǾcJ��.�ʝ�X�����	�k_������G��h�U����j���E�Z�[��ɢ\ز�!�)��a�
�!מ"}ly�Ĩت�N��Ned��%�F��t��#�?A�Yg�v`�l��O�G%q}"u"�n��[2�� i�ТL��!�ܭ���%O�s�F9g�va',ى��κ@ngT���� n�����q�9����.��U?�Z��ǧZ�Ͳ��K[�|	M�e��laKo����?�/�{�U��:so;圁tf������~�����~��}�ض}�[e��˿��s��J�-�����:�ny�z�i_V���ӷ[�uݲ8)��ډj��WAus�ު���K��w��:�&���K_���k������0qx��5t=���'�
��ʅI{١�Q�=Bv��-�����5
�h��>�؀���%�]��Ǒz�=�|0�^N��(8��8��F�yP��A���Lm78������A� �Q	=Jul7�d�������Hhl(6.P��tt���m
 �^�s�q`]�dv���<(6�S;�����D?$:�M8�%`TOK�#t,�F�&"������AC�C�E�6j��	�SB�ȯ�c@6�W��EG��(���CL���Fu��Dǐlʳ��4��rv�/48�˕�C�d�MH��JD��|=��Sv�, 6`�>�
4.P�"c���D"?��k��>��� �lA��p���F���ic�C�k�!Y�:��U�q�j_�02��H>���C�_h����D�ip�&ֲ��t+���K��
x_��n�i���_�� 2�Q	yrce�, 4.� v�h\� v�S�qf�.�#*�*�@cH�C�oW�ŋ�g�ڦ2�ut�Ѳ�>T����f�1����}�q_�zD����6o�뼩V����PK   �l�XN|jo�  �  /   images/07e09445-3584-4801-8c96-91d92a49cf18.png}Wy8�o�� �ؗm,c�>d���5�5�I$K�%K�����wB���ƒDh�ZB�N��5[�^�����}��<�yι�}=<��dan�����X��z�s�qne`�����c�G����g�5��~q�y�/H�.���fP��]($$D���v���?N��g��U~��h���-�tf������x�����W��M��,yR;�{?x"�V��4׋; �Jg��
�����Ҕ�A�d�>���cǚhv��n8:̜�����yx�p�ս=����j�o�������E�"�{e`�;|���b��BJ-�6aM��a�r��s�����	pvf�����^�E���ǯ���$�"���kX�I�	�������GGVRy}�����|����Y��Z&�=���l ��E�ҷ-	k��K�}~7��xo�o��&$���2L2@�C�R �u�hM��rȰ?(����vo���h	���E8u�_D5��2����$T��q�.�Ȋ1�r�${���p3Q����V��a��<�b:ҹ�覟8��/d��'2�=��U�5���b�x!�H������v��Y�^x���N�:,�4`����N����� ����<#LY=�F2��&V���D���|�b�slUO֙W���*D���q�p:Q��*݊�l���-8�Ѯ@��i���;�Zg� ���Ɩ8��O b����b
�t��q$ix�Z�9$�͋��X5sOI�������jd���-u9��%�e�|X��<a/��d�jzz\
YQ�+����7���`z"4�]��ze����]Ñ��lD��.i8<�Z�	�J��W-��"KRc�����@b�W&�i�7ָ���!��	9F��.p�'�h�CцWF�9sQ�l���x�� K��9�:,/��͢6�a�266^j���#Q�e�ě#��.����:'����v�"أ�+}�)�z-z��I+��Z׃q|t}���f��$Z��YV&(%m�}����g�G))�����%h���Y@뿭�Ī�yLn��b���C'	%�_.�8���YYM��]r?��r�N��J�M���"�N�-��?�_sxx�C&�%mll�{k�;j��W%_nT�3s�ϙ�k�q���C�+�·�"uuuά�wn���#Xħۜ�*=�RBP/���Ӏ�)��2���P���N0�޺}��}0�!�Y��k"�=I'�oVǸ<9�(v��ރ�v%^�-V��{�C��m�}�Y��%G���u�)/o~5�ͫ�-�ۉ�+����E�od�z����a�*4�����E61谉�l���}l�׽����whޔ��y�RٹU]7��x;���l(����7��U�§<���#L�:��ʋ��!/��>�a�P���H��V/����z~W5�o���Me�>����u���.��֠���c:{��h:�dd�$�"�d���,�.65-�6�cG�r=gu�śT��L4Ø��p:8��ٿ���Joƴ��Mi��pYu}`A����X�.c���O�v�p6{���q_A�i��دk<�]�W�v��X�.��b��[��o�.�v�������S�}���5Qs�,�:i�y.')��tf��p�q{����C�G�G��v��M)!�BV!������m�b1tȡt��]�6.�m���[���lQ(����c�}��d撾T�WS��/L��ݞn��¾"��>v�tR}��V�y.�7N�1��h����t��l՘e�I��.D�O7U�[~j��D��>�zϲa��m�yZ2�d�w�Y ��Pi���k�Rg���Fǎ�+5�G0��w!s̵�@CT
1�2���W0H�T�%ȓiu�.��~��F'��sr�����1W�Jq�\ϡj^S���P���?6�L�F\W��v�FF����{��U�:���l��/=� S�e0鱴(c�3f^Ro���;��)ٸ��?�V��]�i� ��mY(Flj�1�STU[�.��������V/X9���O�@殉G�b����u��^~�����e���X��R�XRI�Zav���n���,!������,@�kލ�p�S���F�\�v�1����X`U�����oQ��ӷf����y2g��*�[���3ΩY�����'����
"��.�l%!�Z�^x2`�b�r#|S�.S��̌�_�.�>����F0�+�� ����2S�8���rb����K�.~�cw���"B�l��ЍG�3>S���@n�M��M�3�kS>�R���:{�2}Z2�u��Bo� 6�Г�y������{��𓼌&�V��k��w%����@���d=*����Wu9c�ꁑ�Axxg�LL�Ny��[��![��̶��4����!4�r����!q9�z
Jg�ĳ>/z6`�}��m9�k�����˖�NZ���4�y��RC����P�|�*z��X^.��Xf�x(0ֹ�U@]ϒv��?��i���It����L����=���ᴚ��2�Y B�~u
M�lh&�/��4��d/���cƄ_�&��%ڪ\5(-����gU_��ퟕ����Q�	;G-��#�W)��#���/^>�"�}�L*�S��7�]�ϷM�����=�T�)$��@�Y��� ُ���q��,7��c�X�K��~�7����GEc��U߫G��9k��W�nv,�G��9��#z�T��v����*�.�m	"1��u0] <o*c�g�a�ʍy���dI�z��_G�UNe��)�ui��8�82dU<|(e�R�#8��2�Ϟ�/Ї�*1,��-�8ﶕ|Й{�	��ڄg����pm���k�wP�$ġ����!/�X'I.�΂���յi�XX�&��"\����[�c�b}D����Ѿ(�4�v��.f�q[Ľ�D=�\JB��=kh�u�db�Jc֩4�b��r�p���Å�e�>6�+4�v8�[��q?44�n�������H�:)i�+��S�Xy �w���>`T���G�r�k�Q�"�U9��5�)m�\���!��Tb6]�Ϧ�sNJ2�
�=��j#?@�h�s�o?�y�p/X�L�\n�/+���>�d�$��U�m�2#tA�p7�Q[#���W[k9�E%v���y5R��5�w �&�]���&~��h��Y����"�=���e+2�Ei��蘙���s¾���?�T�EcB��Ξ��)}S������ƾ�Ґ]o|D@��X�\�#�N�r`����(\d%���d����E��� ����J��z
�'|kkku��j� �X��/�����mW��Q���"0<v(����8 ����T�!5ﬔ��2"w��䢹^T+��ѝ H�;����>_�Q��gA#�QN>/�
�.w�"㤬)�eb�IK�$bPj��E#���f>�ʫ���j`P�=oǟ��V�&޾sG��	���JH���+��f���n���P�_͚TS�����c�A����N��������e|o�b���Z��Rt4fV	o|��ieOO��"��:�GNpq|<F�I�Am���VV|||���j:�J�W�R3d1R�Ku�����������W��Q�����t��d�U����O��(oIH����jˎg�e �՞�&8���yMU4�I~�Be�
�D�a��a�r�d��u�i�Z����]���Śf��`M,-�=�׳��a�m{���0��V�ؘ#Il��2�ܞ6�#(���jD�d -ZE)��	�l[��;-�OM��Xs�_H�*T���#�kD�����0R�dKć����-�IA��^D�� ڪ�T�`���4g4C�ѻ��k?�3S��0�%Fh[[ۋ�����6ڶO
,�>�f���/BV�a�J��׮�
6&�P�+M�g���'�?p:}�	��%�~���g"?5��|E!����L�|=����P�
Hˍ(�;mpכ��1?��A����_�F!n�hD_����k��0ِGH���Z�h0#;
�_U�������Oovr�	�ȏQw��f�3�H'6O�i*��>0��:�e������χv����^3
K�PK   �|�X=A�'>    /   images/184639ba-f95c-4173-b99b-7b38d7e1948d.png�Y�S�>��hDi�N�;�SJ���>��V�����.�.��FB_�~y��wgvwfw���g���l���.9  ��Bd5�y�Z��gͱ�~�s�� @������ik��y��{h�X{x��[���9�`�V.�6�gb�  �'������خ�qHG|�;p,�~R�f����B��6�=<�8B���b�ŉ��������ʈTl�%=�WF.���R^����N�dppl�c�k����MU'�Lk=p����z8P�]��������
c�XE9"��߻	��1�N���9����u���onS�B��YNK����@uþ��Wl��2�&�V�5��q�T�O�����Ǭ��Ab���W>[��aQ�g;�W��ꎧK�E��cA�.A�	�~�F���o
]�\�(�w�r��7�6����J�UU��My���...'����(��e(��W�]Ե�l���Ht��`��o���{g[��H��;�Aw�w'�C���4�vs4cO�􏯏��k%��A�Ӟ���ӜN��p�z�J/���c��YN~���_<���n��$�?�DѲ��VÈ�����z:e�H�{ÏL�������'�?�(͠��@�z���)��l��j��*�m�뮀C����������l:��~�pѕ~5�����ّ��~v�I��i<fO�a��fZ�a�
���RP�ƴ[�j�����t�ʀqo_r
0�t�)�x�_��k?���f�D��횯Q7o��_���d�������U�F�d�V1g`�hB�+٧J���r�\"��ԇk���Ȧ�"��7�K�="�@�w������|%@�_���[�?�pXK�]MT2��!\3� ����,�r~��|����a4-k��\�=G%��g"°���h�O=��*B��Љ�,�y8�jw�X�c�D�=<-��D��%���jM�|1��|�H����mf���ط岍�-܈?�f�'�I-�F5m�W3yL�/'عh4����K��Q*�Ӱ�P耴�ňZq�S�h]�q�����y���Q�gMnl�H���؞i���4����[Y��6̹O��\@�NRl�VU*Dx$&d��L!WD�w3!�u�\?�*��N�ͽ�T��aѬ��R[/H�(���V!��G��w]����^#����-�F,ol�gkmՉ�0��֖�U����"J1̕Q��J^2q�j��=��z,"D�.g�4�Vx�̣���G�d�t5�T�5X�n�Z�����Vkb|+���U29�a��E�]T8���ӗ�PlO{�g����7�(��P8Iii�LW�&ZH���s�M�U8�Cp�~]o�������u# �{�L1%
a=���eT�k�9��C�Z���=¸�MC������R����
<��[�H-r+�x�",�W�l���?\�aC�X�B�B���]͝��0�pV_ܷ��j%�C�^�X��?���ȟ�̙Τ�m(��il'��0~��Z�(�� �ДKՔ:��$��:0 *R�bd�+�]	?�G���>;#M�<�Y@�{�ۺF�!�&�9.-/;U!(��B�J����9�]wFq�ma:[8F�ƛV��~��
�ר��h�y���*�Ű���ɸ}pt-�m���᪢�#/)a��H�������Ya��2s.�����	��n���)5# TZ�h��Њ�p��UnDѱ"N.���y���{��R)�	�(w�pI��eYX�"�UgYQ��|i�N�����ʫU����DI�@Z��c�Y�u�/�m��<{���g���O1e`iz�\�`��T(����,���a�h�����@��U �auS�U�}ǯo���OV!�����G�yQ<A�\�%��O<�����L��.��L�ᣲ�a�tc���WJ`zX�8~��w�E��W�X��0	��݌H�iQ@\W�@¨�zT�Ūn�2$W� %OjW�����Ls�/�И91�^���7����c���V��u��v�Uz�2Vj��Ξ���r9aP*<SI��;�P�tv�?_��|[����YGHZ$��pH��F}B	�LZ{�-#�o���qp=&yAҸ��z���R����WnA�s�2t���%F(Ja�7�b� ����F�V�R�����
̡�|�D̸ڪZ�ܰBԍ{O�Te�r<�+�h�����J��c��f5C��Y���V���w�oN��|[��8(������1L������Q�83��*�G2�Em�2����Ͻ��WS%��q��ֹ��~��{3^�3R�i��~��,�M�����o6t[�´W���:ݨ���}q� e?]NpD��)j�9;h�L9�Pa��u��d�P��=S�*.��������B:O-�R|��P>Kg���r�c��X�w�����&U�����9�3U�%�%��g���2.��P�W|������ zzs�-X"�O�6��B_��/+��c�]d���-A������q[ �ǥ����J����R۷��+�H	5M	K.yo{V�z;n�Ơt�><J����x���`H��&zz�QU3�!��$�.��g�ү�У�v �c�`�����%ZE�q�R�.;��i2fEH'`W�+�eD�P�����3k���(MDh��D�~�R�B��r5U�&����I	�؄&k#0�*��QWd�n�1Q(���-į���[%�:�`�嵔�]�J��\k���W�^ 0j ׉�%ҷ��n�� ���.�v�rC'i��������Ǻ��9e�R-FY�����r��$�l���d��SF������.̏!����Z��7X�U�����H�GePoN����)Q�O���e�1��L��I�D>�G�#c�2;-�N�5}��P Ԥ�F��뇣ۣ.�����2�4$�+5,nf��4��]p�U�=V0�O�y(�����"px��ח�y�/[�J�՟�"sY�$?������AX�)H_&�;ig*e�ڋ�%&��d%\=[�$��,p�"g�s��h�)k�$�C���r�/��!Q�~�1�$��v:V{�oZ����x�b�'�>ںZ���g(8��g�Z�\�9�m7E��>�V(��D�1`���l�`m�i��id�@�k�n,V�$������Z(+Sp����0�����È��@H Zs��n��k;�6�����Qc�����u�>�i���u�ϳ�6	%���F���}a���`����'�ܐܹ�袀A��,/�ǎ�e�������n�^k1��� ���\��S��֊����[���P}� �9�\�+�$ɨ?��ݖ��9�OvR���P�P0Nh���2��{=ld��1'^|��L?��Mj�N��.�)�&,�9x�+�# ~�б��r��eJ5��~ [�#{BYS�k�r��Hω������V��P�Pa~^݉���z�篪�L�U}����C�_t{���Auvz]~�Dª��c��c�ټ�6�7G�7,���m�A7E_��; �;=�D<p�mWm|ː�S^N�OJ�ˋD�Gr}�+}��ql�h�.W�-�`�ǖηչȖÞ.\eD����jZt�"{0�GA�w����4d���w�\�pD��n�mc(�^!������?����T���35նn�[�}���>�ՍeaL����,��|$ž�(��22T����К��&���Jc�	Ҳ�uT�b��0���� ��:��65&�	(�D�|��:�<H������!����kƝ�7i4* ֶ ��E+)�_�*����T�DJ[�k#85$�RD�|i��O����^<��&��{YgҞƘt�9��T�&j��f�7���(�0mV�6�.�GD�'���T!����
7frPZ{���d��1��Mq�lϡT�6Q9'FO���=4�"� �u�e�¾g�R>�T�2���X��n��5��"F�sf�h��?IW�ȷ)�L�>�z��Y��F霂��zC��N[�O��oG-Z0J`ak�Y:���{�Ў��f�&��q��m&.��Ǆ��e���j��#�I��$�/�!��X_�ﴆ1�� g0b��"�V�����RR�F�o�R��{��#-E*LH��5��"��S/�ŀ~�
�L�D~�lrQ�4����	�j��§#��,����-��h/Y�WZ��NB��i�O+��FB,@-�/�u5O1�7.Z�:"t7@�Kz�ONº)��F훡-`����΅�����G� Dg�.�,!fHW�&S��EqPB�֘��)��9�y嫆ͅg���Ao[��'|%���;ʰf@"Kx�HG�O-ƣ]��6����1I����HR�ETj�y-��$!����W��cuh|��Xp�}xn�_�������M}���*=��jX��L�%��s7Y�*��:?=|�6�qW�h�4��9	
��p�J��0lmC����q�0,i�lɾ?�w��Q{.��&K��&/���־�O�ӊ�z>�}�s\u�0&�㔢7g�w��`�ȸ����݌f$l�E<Lew����/�ց��M���k3�9�K�υ��,Z�����ʈ�g�c�@~�^�D��B��V_WPQ��Pe�I|�k��R� �/�RD��<s܈T���J���ʷ[�)���y�eǕP�X��Eݕ�6�V�unC4��ș���k�p@R/iq���ȣ�i'��q/��vp�H�kyڏY�][Fu�j<L�8
���eQ��c�*��CK�N��uy� ꙴ�G2��������9�liF�
��E��E���˔2�q #���"W���TX�ک�+9��n����
 ���>S5�s�j�S�K�Ff�q`U�>C'z�6�9:>��W�L�m�8�1�:����]��l�F�T�7�g^����h�KE"��U����CȊ'W�~W���l�ă��F�i2��PVpİ\�� ���]��'�FϋI�7��v�v)f�IQ F
�n�{ރ�� ���(��3��)̹�v�ľ��a߸�����?ǓŞl9��b "3=�^��}t��ۗ�����^I����5�)k��E���[���%��~"!0�������*�fP��*)s�*M���\�rr���|�(dn8|��p�mɒ�/2A�r,샢�kR�i�?7��/�4vd��%�w�yR���`��S. q�	�+��)�5�/����.�B�cC���f\���QТFɽɱ�����/���r�yzA9��h��1+|.��v��j� ��j�+��;�0S�TRQ�e��>���r�G8,��=�����0$���6���n�'�L�6@�X��Y)K�8��C�۹��ba��B���h��m:�C�H�9�q�,���K#I���(�0�wru�kA|�~��|�H�ȋ/��_�i�a�<�QG�R�'*d�r��l���s4�x���9X�;�M1������Y���F�\y���֦#�܃_��fg�p$`���,`ӧD�����(m�F5���]A)h`���X�r~�2��[ʈ_8]Ѿ��ya�TwO.91·��.��r�pf�V�Hvm�G[#[�O�x�v\�b� �pt4|z`^w¤��u���?<��G+/'�CȚ��r�hLoZ��;�(xK��e�>)��n�b�������D�Q7�
	������Kf�3O]ض�[kh-
�5ޝ.�@tC�P�m5W����M��|W)q����R�ƸU�����Z?�vg��R^;�?��P�-���I�+'700b��^�-x�MrQ�Ȋ18�%)�^�5D�c�H�S@���]:�����Z���1�8��W�dQ�R+iή��QU*��,s���0��WRN�P!dzײ[PG�i��U1mvI���9�8)Ɍ�w�j~����66���s�	q7��}
�����K�E�5��j)fC'$�c�y�TC�h�|�g�u/��}i�����.7�3��u����1���/N�ܕ
~*��ԛ����:��-<�!Z�Ab$ ]��vU{`�}��t��<v5�2�`�{�8����|]H��o��\r�➮^
��B�|�.z��3C��RY4��� ����$���+e�����Ri��wV�i@�.�x[{�@�C,�1��H�X_=[TE��6��8^���۶�8����,ˆ{���>~�R����~���0�"���VO�2
�a�??J<mm��t>f�@32��uS�+�@�t��q�2��ux�osލm��q��2|�����X�Z�����5%�"
ߧ3p����d}�b]��n�%4�1	�A����C]�㵚�b�0��Vv_����!=, �xyX��h��`��6�&O��NHj<����?���D�u����溴c�>oM�t.���x z����t��<��Sk��c��;J���O]gʛ�ڞ@��'''��E^��b� :!�4�D�L;?��M���g��-W����I:H�ׄ�����9�Y]m;T��s���s��N�Lח��o��׽����~�}��n_���t���2r���b��As��luI��M�s�������Л��_��m�w%7Ø僯DJ$"���)��.5s�]7,<ܪ_�o>,4s�_��[�
Ӱ�x���4�x�^*��\�}�1���5�tTYE�z{DjW�x�M�aa��'�  (x�a'��ĺ]�P����_�n�L��:2���4��S^���l{z�-�Wn���Mx��H���r�Ϡ����qmCɍ��fԦ���px�ud������ʣX�4+�ti�#��9��ڷ���k �|�%�3u���k���GܵG̋=L��(+	��H̪�_����rS�����q��Q4r���x~�Qz�1�W�z"{��:^� �O�r��U�f��PK   �|�X�wM�|  w  /   images/5e95862a-04ad-4971-a9d5-8bbbb67b4e45.pngw��PNG

   IHDR   d   #   b���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��[	x\�u�ߛ}�ѮI�dɖ��`V/P�[ K)	)I��Y��Y��Ҧ�YIB�HB�J��	`�w[�$K��5��43�}=��b���6���~ߓfλ�{��ι���b��Cŏ��u�(���*�X0�0�U�����,A2���V���(,$K� ���N-��2
ϩ��%d�=3գ�͑����d�O�a$�D���z$4JȒ�H6/�v�$S�,<G�CZY�,����d:!S�L2��Q�A2���d`T)e�0�4H��4�j���zZ��Y(Y0�oO��=��꜐�z���X唸��\X�/��%��g5�\X6M����@������.=>�J�y����(#Z�i|q�e��h��֌��۸�^��҈NM�o\�@,��ARc����.A,��w"��"�&�J(�����ï��I��K�C�R�;{݈�m��N�߯^
�^�o�я0�fS������l$Y/���}�-p�-����pǵ����KW/��r~qd }1F}^�eZk*���=��!�'.i��Z<��	C5Nz���R����ڏ!������l�bC�<���B�2)��dƖ�Mx�@7G�4����V3Z��ў�8�1"��8�=�J�!��St]6 :�v��3�^��v%�ռ�Յ��4VV����q$��m����-5��=�Cg8�;UaQ���^����4nn���T*	�� �����m�z�h�l&�~�-qر�n�T��Ƌ>kL)e!����������8.kl$�7�l�[L�xES�t�q������t���Pi���8����26.n��V$����XbW���4��ē�i4[ո�m14Z�$�G{è7�غ��,߂�WF��� *�9ܼ|	1���Z��Ó�Gx׊�0��}uf:|4�tX�|	�r�Z�϶� ��!��}S��w�������е�.�$��t��֔q�2�h��߃K\Ud!A���xv`�x���s��"��prW6�#���i�r�4�"N�t��9������~��EDe�+�06�A�Q�l�)̹(�B��q�:d��78(,䩞	�H�JG�g` .���`�x#��+n7�*������\*�����Bv�M@kv�x$�]������w#+������O�7F�d���^\���:��j�f���_Xȶ#n��τ�⨰��ð��i"1�|�3�L2!|�l��ڮ���E���w�x���#���RTP﹉Z����/HFMIc����'�"M��T��+����_"���D�w���%��dw=}X���d)(�g�W���4�>�Im+y_C2�dz�K��+�D�>��8���@6�g�g���}%R�}�e7��QE��~�$|����CN�gͺ4b�Nd͸���Mu`&�>��h���(��Q.���q|�Иx���g��C����Ǎ�	��q�u5U��\>d��1���i�}�d*!�H9(Ɋ�s�XQ&�j3.@|�sd�/q��O �Y�dL�'�̑��	s�,M���j��e���%!�jRĘB���X�S$�䌹�D9h�,��V�K��O�K$�>O�g�p ��頣�ٍ�����^�ɀ@"E��ra��Hg�qs�y�u1y!c�z�)��8bAa �d��{kG����G��N�)#�����W�⡑P����k�S�(�=؋\,�/_��,&'�����S�㮚�*Tu�~Pb�,>��ax"	5�d��&���s�x���t�|gu9�&'�W���4���_�34k�ZH��i��Ql2�1o�ef|���J)|��q��M���j����$�z���U�p�f8�,��he��b����`��./�$7gIl���[��9�ܝ;w�w���iTJ͞����hr�׬Fc��~�/��ؚc�OR�7������'{:D�8�1��J>��/
Q�c���xVlB�h�����)Τ��J�@Mõ�(	�/�h����j��_�.�M���j�9�����p���)"�IG��MMA���TUE�e�T_e���*��#Bg�{����8��R��	ᖟ=����J.�M�!���X�gs$�q�Ex��[�l�I���.,wV`��<���׍�>|ʉ#&�>t�*�<�Οl�<}�`��9�ʁ�BΎݘXu������G��rĳ���А�4R���f21�9�M�&�ڟ��3t��ͅ�\��e�������8�����KV��������ɬ�q>���ǅũ�m۶E�RE�L�4�\e��z{*��\��N�2��#�reF�"� #N�<N3�D��_7]�o�>���y]�+������nć�Z���Y���_a��Z��}�}�y�
<��4Ƙ��<�E���f���EL�$PL��E)ؾT����'f�{؏Z�hB�(Զ	
Vr�)Yh(O�?{��i�q�)A�(���:����M�N��r�l&��?��Xk?��*U�-��ɩs�` ���Z���܎dm�2~�/o�(�Q7�K�� ~��q���M?�!��L*�A���qw�[��/_��c>|�_�#��~��uƓXPf�/��J�J[��SG��=��aQ ���8�Wfa�,�F�pv�>oP�j>�܉F�_?8�@2-�g���?FYug�����Pj��C!�l@<��ѩ0C͒$&��2��P	AUy=���$v �߇�+�K�Ť|�+p������@���2
�$�(�]�*Y-�4��y��ب��*I΅��*vN+���]�oN�)� 7�5�gn[ۊ/}}c�~��Ø�'E�Q
��]X�eF�`̽/@aKa���ܠH0G��Q���w�=�w �kO#��a0G�рϽ�@$�P0I̹�6Gt����;��^+!G�� #,�r��:�g�����wj2)�׋C�(Q#4�L���Z�
v�]|PC:r̢Pc�p��ۅ��w���phԋ%�e�ޭ�1��G�Gﺁ2g~��Q�s|�F������u�NS?ʆ:Pq��`� %6��)l)�s��yB�c]�13��$=���XPU��lF�e����0=�9g��ep::�Ik�tRtf��W1���5(�,^tT��)�)�&''�u�V�V[��A�T$�s$g�T��]��?!P�p���N�2�Qr��Wn���U�z^��Gv�s|J �N�̉��\�(Y�!(���8����H���
��fG�Uyx� 9UG0M�n�z��~���8973s|��.��%��{Ӎ[�ۿ�`P���ɒ?���z8���1�E�|����<�BQ�:�|LY��s�x���B����m6�#r�$�E��?H��尰�@4���%Mjq��õ�ކ�
�)ُ$��nh4��E2>���M��,QA�A��!����[J���
7�m<�/�+�&�b�(�� [���i	��^��������&������6�GF����\�K��[��+�yi�Cbu�%� e.�N �\>>��_P#P�p��S��J@��"8�H�$����/�=F�,mh�]��b64��=G1�R�.��A� C>o0N%T��MJ�i�#��>�x9���u��o�X�n_�䔇=^���| ĺ"_\�ڊ��q
TLU4�9�U
	1��@������?�[�uq�:��)g�|�QOɑI(�̤���.��)B����)��&C�Rg�oN�0�,QS�e%�]�i�L����A�jT�P0�%O_ATck��l�N��X��
��Ǐ�^8��6�rڑ���4	8j3��}"Ke�P
�SLl����n
��I{����âH�����d!iB_��[@�.���:�	��L��=-dZ�Ad�0�q��e�4,�}��pq�;�4ft&L7_J���,�+g��7��c3D���(i�ry@xIi�f}n�kG�X`3���x��}'0M���U�E�R�.��"�q�_���T/�Ȕ�#\���'6�������
�P��?���/B46�t��7S�HE1N3�PX����[�^t�>�%�J.�0Y�+6�NH�̼���8�{\���j�M����g��r��3�C^f�%|���.�N�^���x��$Y�e f(n޾};<6n�H�Z>2hkk��l�� 97H��X�|���n�#wn��f�Z��w�`y༠��ږz�u�B�A|2<��C3�҂�(&��[|���x��|A9�faig��v��e-��L�l[�HT���T
����۪�q��n�:�N��qK9�떣n��H@0E����µ�jt��(9!���EMM��̖��-����T���䬁����*KtPO�ܪ��W�{���������c:��f!�#�ѓ%��[/}A��[�<ϒ}�����W�H��I�*y�2�Ǹ��`�>Ӌ����f�)����saE��k�N����-��73
=%��h��Se���ǡKF`�$�f��H�a�;������9Y�Y�U���aӦM��gf�\*+*��+ª�����rg��^?z&gp}��Hvx�d�/�{��&����G�d9q��h((�R����v
�G�9���
G���&.��n�,Fa�� � 7�[��X����T�2�ӄ�%N<�l��0~[m�������fo_jS]QQ���Pf�`�b_�E�l&+eiPY�%4�d�D!Ic'?rZ���"������r�����������#�QԹG] e��"/.�	
2�3�%܏l��%a�=���iIRUؑ����84�Ǜ�K~U��xӔ�sR�ۭ\o�C08�t&[b .�H$���p��Ϥ����G��t���qU&U~XSi��tj���i�V�Nf3��%������s�#���X��4���E�"(y0L"3Oث�	��&��̊0M��p��2�Ȫ2�h~�B�:��$T�v0�$�,)����l8E� ���!�I�9CWjr��n7��,��1�
I��~�UqlD�����4^�Ib�7~�Q��7!�/%P.N�׷�d�&���^�5��Օ6�8�{������W���LY�f#J��$|�t�o!�lSV�����v��]#����Ms�bC�?G)�¹�D�-��F�HȒ��S��v��
+�=�ª��weeqd�7˃C2�]_p�Q�����ZL�B����馛ć9GI���aaPhT�Mk�[���|`�T���SYx����h(�j����Tr�b��du���N]�ӻ�5z�j#��L�i��_�_��%�e�����=(��V됩�G63KX���r�/<��-[��H^o<�fE��g���Ô��]C�����D���3��g/�$Wȶ����E��\������l2��Yq��M2%��Y����+��:M��{��~0��Ǖ��8���b*pJ��OW5;�;6�[_�*&�}��i���0�lÂ��#AH��v'�\+�0ցD8@�b)�������y�/�N����bO����ɜ�r�M��iY�R|B���MG���I	H��h�$�`���}q��2=����j(r��'���bT�K*��?��D�8�卦|T��f(�~׋�jq��VNćsj��L�S�$`R��a��*�����:�}�W ��~�,�H!n�zljva�|�p0�N���rT�5b�)��Xі�qP�x���ȟ�}]W��6��5�tOC��qe�
�m\��@;��p�2�����.�vG�M��T����"�H������ِM�˛W�ŵ���,���V	e|���9�{����(5�z{?R�2�LO���`1���>�)��iE�Ռ��9����>|l}�8v���.8�V����6cYM���1ʽ�~�/���Y��wã���O��8�����w!c�E��>��W,j�O�� �qIl�T`����z=�s6M���-f�ж??xSj#��(>��
��X����PΎ��Y���4�����Zw��￠��"ܑ?����.4V���v�'q��Z�0\hq��8��Sqܱ����huQB��6w75UbIm�8��5ƫ��7��͵�I���.O�XY�(Nd�����4���a��Eb[���Yl��*�뚚I��֖ v�e��ʀ+�[H��{�B�I��
+�Z� �l���865��	w�\ �V4����TGq��VR��<��a�Yƍ˖�̄;W'�.?\ௗ�B���=+���Z��]��`4�q��홁d���\���]��CG<���W��a��kd��k���d��5�����[�~oG��!����>Zki&Np���w��XU���l/([���1�_�7�s'���uxap�4O D	�S�^��j"�64�	�yf`
#q
���;��96���^u[F���j�d��To
q�n~�5�#�\�,���j���1���}�w��>�7� QN4��o�G�F��o�L1���}X����84���'�W78��'�M葈����=��b�7)ag��4�Γ�!z��kg�	��R������<��k 7����(j�8$�V��L:6���QV����E�8�>�ā'�ů��J8�	����7�E$�G��m��O���j/�Y����_P�������~��*>��C/����qX��h����랝GE���������;艄�����(�t���?_>�?��[�꿙���� �7���?�aP�1��Ž�����߃$S�Q��o�iߐ��Q�RY|y�:8�@&N��W�����D�D�Ar��:����<�M����E���j�_��,�0XQ}os    IEND�B`�PK   �|�X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   �|�X��O*�� ~� /   images/bd13d416-9901-4cb8-93ec-096849d17163.png�eP_�.8��k���� ���58�]���www	�A��	n�ߺ[�[��q�m�jz�t�מ�yzz�����a(��U��Z@ ��Ȉ���'3l�<DZA�|��#��(N�u! e��L�gu`'���������З/_�?;�B�L�,�]�2�EIA *�����G��Ɨd���(n����v:���V!�olfdk�&pCp2�Ĉ�P�_!͛����<��&�a�0���f1\S�qQ�*Y����VeM?��Q,hn,�=�G/0�8^��j��o��~�n�9��D��H�Q8�?��#�o=�_h�s+�aub��w�3�ϓP��I��L��~�������_�6I�1���4F��h[M�"���W�B���zo5������|v<��l�f5�&J���*�8���q����|�*���/�~��nT��uM3��������C����h,������]�:���nZG��W,s��W���x���������;��X�f׭`}��#��R���	�=)��粲���g���Zg� ��٣wX�/��Zƿ�M��n�ذ�9�����n�h��]U��0����!�G`��۴z�v���:�+%�*�r����߈��"Ø���q4��=�?��
���O�Kci�$<O[�d�l{�/Z��2����2�2t��3^'�?6�l������4m�ෟ�s��4�'������?���ra!#�x�|���ᠶG!E��B8Q<������i��(�1��4��?Vp�D�4���Y}���#���b �%�94��`����T[T։x<q~�l����k<�i訇�jƴօ|0��IJ�Zy'�A��T�2X�ubL��v���i#G����Y9N��ѭ���9��cȈ��$�LA0Ȉ?=q�L',"8:�GW�|L����������/�R��ڢ���w�&H�+\1��3R(mP:N�0�ki�3�R��"@�&���d^'K�)��wG�G^T�J2sP�E�%r'�h2�!�J:촳$%p��&0tգzKz�7��*~����a����B�wq��|E�
;�h��_�>�	���Jz�t�#\vX�Խ7�6M72׈4矓�s�Gj��� "F�t�ߧ����O��R���c��P�Ӷ��P���g��E��j;�,5B{\CuR�@q&��� fV0l<�>��2�%04n
5�-�	Z\�������tu�]Ł	B�����P3!�ޘ��� 㩐����^ڽي�O�F7�${����Q~lg���U�{c�x>ǎ~}�Rȫmi��z�����r@vB��ۄ��;K����0J�`B>�ꬰ_Ɂ�+8��X�T黛øQ����bZ��&�?D�>�O��p�ڙ(#0<�3N���c�$Z����L*e��cXLUg�,bIN���G7�w-�%����,`
c���+9L�{�δR(����~�A��)�� ���64�c=8�Q��Q$�M�%�/z��`�U��-f�iK*Yr�0 (�B2=����_n�5o����r�
4�:T|�W�"Z�e$�\pt��~2#֡��3��!�U�7T&��7eOM�����H���G��6qL�%�QWVDWG���
l���e�kkS�^o��E����R�gjI簠��9�/�1��ף�j�Jfr��ŋj�N�N��@Һ�4F#n�h��vɆ�_ڃt�\l��AOW+qt��k��0�/{��Z�:Qv`5�XmJ�J�"Ja����B?��-_�U@Ȼ� �H�^�ћ�'n����8<���vZ�"r��Ek�r����_J���LL�L?>wS��
&�;s�J�Su�7�� My�k;�z+H���=YtL|V�)�l�̧[WÁ��$&
\����6|d���j��b)JC�BZ�`��r�����$'��mٟ1��DK��.Y�G � K�PD��$�K&׳ � 'Yf}8L��8H�Ǿ?�G��O��n|��z�cZ�2tUH &�0A| �E'�s�S@?�G7S5��P�ds��W_�=R7�27�����@1�n�^��j ���#Y���M�;ic�iX��>��;Vm��q�*��͵ȕ�Ɛ�8_x^p�^�|41
jF�V�� 8�ژ��CUeS6FE*rIrv́H��k,T��bQc���V� �T�w#���m	wB'Epm����d����]��mG�Cd+nW*	`<&F��h �3=r6��B��V� �Ԭ@��j+t�ʯ2��)?=���g���u�l�e�C����t�`��$��#C<M}��[d[�х�eMU�z�BҔ�y��x'#Z��ͪ��K;I4&�>�1�) XL�g����F�k��WEJ3A��"D����Vݵ6T�@衳�N��)�f��$������#��
�&c�b��$L��
"��\EP���BTW����E=2�P��l��d.'���R}�e�2X�b���]�u�9�/�������U#V���v�51X~�������&�V5>�7ԝ�N�p�Ǯ^�L�8|���y�U�x?I��g�=M�-PDs�Uz	�z*�}��M�4˖q���|��[/��[�-���D������xj����/��Z{����}���m[>|��Wӏ荢0�Z���&U�3�C�Y�OR2&vnK��I�H� x��>��LOm!	�6����F7U.ϊ��e�lJ}׾w��o�M�}��A�����{g�tR��C��y�i��b��|ɪ5��i��v� 6��� �H�(��J�����Rq G��:�q��_��z�XU6k�����M}>�D��.��,�dH�K$��ծ�e�Ԕ2��ˮ9d�����̜��K������	�R8Z&�71������nm�N�}�P����Q�7ٕ��KSu�r��B�[w�\�7�ba5�I�2��0�Z�K	2 Q�j6u�����M�[�D�EU��"��N���I�������W>���|Ӫ��5��+W<1� �Ҁ��6�G�� ]m+	����-Ǳ{'�k���EVHOܺO�5�b�t	�dЯw����g{U}v��iv�ڪ����\���:��.@vt`Z% ,����,��6���zk�I���u&[�UҪ����SE�~F�ܕ��(vg�3h�^����͉Tm�:�*t�Qp�e��vp�*mM�<D�h�BL�/n�IN��Mʅ�
���4��(�L:Rk�#�飉v�N�*+k=\�i���b.�J��$���O3Y8��,ͤ,^���9�N����5������36n
*����k%�C��ȵ������cK��X[z*��Z���T��N�Kƌ��Z��u�`p����j�֬��YB\W�⧭l&��p����¿M�[Ԏ��+�+�}NsT�%ftp��1��]�ف��B3���l��ks�P�ת��8��U��k>p��.á���Wd���:�D�eKj�!O�02��gipﲲ:|mՒZ6	���P[�: ��_�ÝM�L����?M�[8w����%X8�	���N܊?��v�;��9Q���F8�.��b���}��V�e�?��	�4F�9��n�*�",k d(ȋfK	�v��(��-��,Jg&���v��q�@B]�7c�/�3�9����_��}��Bp_y� ��f����^4}�y�2���v�5�gˆP�>E�`�nQC"���#����Cu�������\񶕡���X¹?���X�y��i�kp��/P���d2�J���a�z��vND�,�y�𻙲y��r݉]a jW�����jU�H�PWk�%��� �@�2'T��9��Dg��'�-:�ɪm�>WV��?L<�(A]bH ������}���9�.a8��wJ��"Z���aQC�D�g�f\�@}����V�X���,fS���d��M?��T[fO?-d�kג7�R#G�� �o��^�-\h ��ֶ�ڄh3BX��l~�'�3ʮ���f&=T�Jq�A���d�='�� #���`���:%�u�7�쏌����s ����X�1�^Ҙ(���!�a�a�ɀ����=؅pim�)�=�N,#���0�G=�O���b��
u�݂}+� �~�-r��Fn�����#z�^��6^��df��pj74�ű��5_r�O�8#F84��uzA�W����r	T�g����g�� ���a;�u-+\Aw�8n[j�v�������s�6��P�����tg$a������S������p^beG��zL:��� |�:��T��ڂ�����3��9�P��כ��g$���7�(���z�;n��wz��8�����K�dZ��(R��I�#e��V�$7�!���*��<9�73�U��ϝl�ف:���{�b�A�7���Lٵ2aJ�,�BV�ӂ8������6�����Ԛ2����[������ģ��5'�`3V5�n�נu���Ŕ9��;|�|�Ɍ̏G!(𵩦��lg�k*Y _�fr��p�ƿL�*����c$�����S�y���\��<���!Xۈ��~|�]i�����h��k�@��bt�x�,(�
~h8D����G�D�P�����(����pI�����?���.�X�E���->[9�L6>�C4�kh��X�Y&�ګ�?x���@+�Ɲ�0+�h����S>��_�uL�k�Jȃ}������b��fm�q�S_�;�'޷Ȓ�kq��ն�o:/Pc���/�ת)�F�gP��Q�)���q��j�A��M�UMq���p��˸Y���Z�b�V�����&�x���mTT�RYr��@J���K/z����Ͳ�/�K�M�ZO��ߕ�X;o������R���08��4E6�5 �����@�r'�+�0�U�y�
�uˊx��=5#%d��H�1 V��n��
{�J�fV��g�`J����i���M��|�2��P��p��m��W��� ��(�-;B�Q�*�oQd'i�lG���k6�$6�Z4�"���K����m�yoO��im<[�N 2�,Lb�$:�(��h�?���U�G�DE��t}� ѓ� q�N-��@�mq�:� P	5�\���;M��`1�q����_����Xn���N��ؖd��O֡j��<�9A�y �C
�~19I!��%�1��:I�:S�:S�:U��:VjS�Fo�r�*�cw�+�c��j�`!�B�
����~�(��1�ie�-F��]q[? �ۡ�|�tkLNS�G;D'	����
�oϦ��㠟6śƛ�*������$J'1qi��|�ʉ/��Ec�9����LF���w�%�[P�:nov��8{�*>u��lHd>JX���p�,f��.(,��-�qA?n�0U<Z� 7�ݰ�Z���e��A�_��Qiu�ҩ`G��C=ē��s+GV�n^�|�$��F��_*d(�.��>V��+�N�ZUV5�\�
C�xa�d����O����[~�ыE�������҆��p��F?GC�L�uCYG����X^=<��C��=��y�o����P��A3e�]$rJq#�)c��q���3OB_)�· ��fڻN�l�)��[Z���0�\Q�M�//�0o�TK��fG�Nk�R� *�LemQ( �֏ȇ�q��_�2ں�^޶Wgg.���-1�:��(7	^��p�R�%[���9
4�<�J$�*�$t)7m
�WR ̭���:�-�寱�<y�kӨT����E�Ǜ!H8�Y񇇧�l8�:rp��'����K�zZS�_i�P}Kf@�{��4���j؛6n�`ki/t��~���3��/�ؓF�G	�cE��ѹ�����[�S�)��l� HPܾ�����ﬢD��*�2}UF��������6N����t�'�xrY�l@����n�.�ݚ�i儝~�o~y�Q��=�KG�R>)��onDFXb#�-�;�C<f�E\�����\��,��2������%�Y�}���G�����,vt5)���h�v�r<��7�Ų7�^&��O�
s����P������S`~y;A��[OѶ��Y/��&���L��M�����,3�+��~��|X��:Z�8��$�lq%҆O��g�؜E���������Q0��X���F�e@�%Qɜ�>��h�˙s+P˾-�	�����C������C��GY�,��f�3?R%#S��.˾Y��m5�*�F�f���%��L�Z�h��*��φ�* �<XC<�с�J��KDj�8g��In�.n���͐ǘ��J�N�ZFśw����0��x���Q �����Q�4�\��u��{����D���`�����'��+��j����x�54�E�A�o�Q�MX���)s��f���0x��Y�GNT8�9��vo�r�m?'��?]A6�J�~��N��n4M����k5"&�D|A0��̤�u~ZNt3-Q	H^���c�6N�� �����[�D�E_��@���+[��QM���J%8�h*�@vq ���Ӏ������Cסi,�:��XoyW�{��F
����	<1�XH�ZOv���S�{�I���3�M^[N�2<"y�3�H��&ꉅ��|��A&T�oމ�E������e�҈w������#�n����8AZ��e�͛;��:yf|���fPd�p���٧=h1��N�&������"� ��	z�%vq;f���Lm�e
��z7?�{���' ?�0��i�|�$��/Y�������旫���6좪�U���7d��s�w�F��9��n�h6��p��\�W�H�t�kߛ���(rpC���Y
�tfچf#�_���G���|��|�����*峇���^��7�[>r/���02G�Vy�d�Ğ��r�9�D�D��R�	�v�EǵN�q-YB�%Hn�0�5���B�3!�>Le*Ӳ9���'w��]�B����͘Ԥ�D��x�c���9X�c�'׉��e|��FA�CԾ�zo]-�B��5A���$��:�\:�#�Y�+3ןN�xcZ·��#���߇g��z_rg������,�]A�ɪB�9{)^��DmH�ZlMc�ku���1�+Ē�+�W�Vn����A��	3�ߔ���l�+��YJ�d���КfK�C�<���y����Ȣwbr:f�qz
��,�~�8"��FQHt��Qd�P����FPT�F�8�t��X4�� Ȼ؎M?�?���>��'��kƟ�� <a�6�q
�k��1Eq~/�զ���r:�C��g�&��Q��C�l�139ut!�J��^g5��2rp��ò�m}:�T��/�M.[_�E��X�U��eI,d|B�ɩ0nn�ܺ�.�q]Ƃ(B������_���	?�-Qt��;��7��/�[N�]ߦ�I)z.gH\s�B�t��2��� �5'�0�u�&�����'���
>sF��qe�[w��ss�ѓ"����ϫ{���%���=��`���=��q$�@=��o��KM�Vh+:�7KQD�����	��X)o0��&�?\�D�F��ʩ_DĶN��U�<k}���Ez:$���Ƶ3ڧ�#�|*y��Ӄ��ϱρ~�| ��v���>�;2MV�e�([�jl�:>Ģ^9$�(9g���Go4^�GLq>8��X��^�9���\�n���*"W���4��	a\�X����dsC�z �)�B`�&VI�ɘ�nL��[A��V�w㠻�w���;���YPC�3=r,/D�zI�Y�K�U�/�6h��R!�5+�5">���� by��+*���Co��^�{�w��J[��¨@�iR��E�Y3�3����[��*�k��S�e�Ńn�b?I�w,�_�)_@��������*�C�����c^&&��X��@���'��kr:{�u? ��k���8*Vx�yt�D��?z.T�L�{<�7�m�~�+y�.�q��UJ��W�@���]�Q\K ��:fW�,����{n0�N9P�t�������s:���D��6�2U�A��Z2��HA������,�r��c�_�Q�G��:�mNt�����p:"��}^�;{��Jv3->Dn�T�N�~��r��z���I��m�y-2�^�#t�A�z��ɳ�_�/n�x�G�ƶIo^���h���e{���;����,���,4m'�.�1�����;���hN�����9��Ai ���/�onəڭ]S2z.�� U���.�F�В+I4X��A=����6x|����_��z�7ך6��ƥ_���I����Jf|��Vb�م�?>��t��{!�};�V�,�w�7k8Ń9��j��Ȥ�3���+:��d��@�#xs��ڂ��g8@��}��ut��"<׏PM���ޠ/�nwE��<�Xa{�s�Z��������c��A32d�%��&��/�ŝ�$o�.?yMS��ip�L񮄲+��)C&�]�N!T`&���۸N5��&m�|2�'y)�+3{P�pS�	������f�HŃ>><xC+�|�����z诜��i̜�ןO��p5a�����?t�޹a/$�HF܈�\���@��1D�R�����	`	g�
5;������~G�n��_4�H��K���q/ѥiq�/Y,�ϯ����L��F���:�~��C	�V��PM��8�Pp����� ��qX�[���u#�dt��P^����>'��}:ܡ�5�K�o��aw���Bݶ�Ɩ����6I���{"�	������l��[o���O�-�,�+�ir|�d�!�Upm�|'n�s����$�IߐI~\2q�^�֨��^A�Ub&ށc����ں����i{4W&8������&yO��e�hn�(���i��^��;l�uc��Sۉ���nN-��תij�E�k�v���,��z��o�;�&�t�=����Էx�%�i(��
٩%c��"dnV!�����=_g�?{��ֿ�q�'{~�HSns@N4�����w`�y����}����_�3�e�	t��O���,��F���P�'���5E��~1 ���I#E"�C�2٭������Be(Ìx�� 8�X�� ����%w����¤=]ę�Z�ȀA�K��cU@�p���p큖f��5`�\bɗ�����J� d��(H��}��+���a�X�y�s�R�a0xS��Dx��W9GO���K�>[�hZ5K�������ٷ�9�1�4_z��Z�����v��:C���&����E�6]翣�"�fv��0�_xcێ3�k���Q\"
[�� ��ķ�?��B��r�#\�:D�i8vfA������HIz(��u���u�G n}P�	/��Ѱj�Ap�������=񁱘�ߠL�+��F�I#��ըꏣK	/G6^���*#��{�>r�����G��T�.xӚ���*��A���%Cm���a
Vχ�('/�m����sx�?y1��5X��%x��As��v-%����ɞ�h�	i^.��Hv�9���Ҕj�X�ʙ�Z�tZ��Bֱ��{�+��u�_U��:O�7��eE;��Θ�!�ZL���u�u�s?f�{��*��IB�k�̃$�����Җ��s,&��w����Ө����̎��]#�k��5�n��F�D����,�<�IL_�@w�7��ѡ�mU���6��dGr@��Ssz������N��q˼Ҿ���s�������"���G�-�R�5�(��[�%�I�U�x#}��6/�0	d�lcl�6��Jm��\�fP��J�6m��'�<x���1��yZ�PE���?, �M�
���`F[�v�)��6O����z)N�6���7I{̐�vg}���T=�z��{�D��>�����+;)�B���
9䤰�n��؋�jMW,)�����?�
cG�l��.9C6�p�:�����Q����������˱��p��5�on���ʮ2���'�/��N��͘=�Za�E#�f�Y�u�c~��X�U�:��<ݙi����e�V�ԏ\��E7���1���On��u7����n�}s�󇡂�ߺ<�ӘOk��OF�K.����$L��Mm%uu%�c̻��7�h/	��X' Wr�<Eji����:}0��Π���O���o���&K���`$z�ӑ��ZQ��y�Cb�ǔ�;|8n�� ��g�'��΁Q)1Hr�k��>(_���8�/��� �	�[8Nlr���p#V�>돊�_�N�&�����߶�2��ņ�8Y��qr�>�OՋo�"y�m��R[��N�fW.���=Y����]<Y�P�jMah"����A��}��s�K%�1�H(�p	 y�7�ZYw�\������~	����h:��fO���$"�r
�G�S��-A;@wboӯbQq���A�P���
�B��� @f����-��/��1���nsJԅ��*�Ŕ|bQ�tJ�K�GF$U��R�����nE���CP�u�$t���%����H��Fr{o���ʽ�~��!�x���bV��p�JcI�ؚ�p�}hk���%����P?k%>V��Í~Ш�Ø�ܮ6)��GI��F�:�k�><�����M�ٍ�s���c��;S�G�GE�Ɂ��R�t�I2j����M��
��$K���m��/W+�ԑ<�Cj�}Ύ����)�iԟߣL�����b9�c�[�qf�-_3%¬_��+�4HPE �N��0E�֯�k5��lm��a��B�Δ=��!Bwm��I���}y�x+9+͵���-a1�M�D��^#a�E�:V��[��V�+N�7�hqaછ4��+ǷnՈ�~�F��ŀs�7�+��@��L��g2IbI:л�px��&��Ѿ�mv�	���X��<%��n���%O�5��� yx�� �yM���E���2�?�����<��mU�_yR��V���v�I���|�sA��м�����D������.�xIz��c4W�*u�D��z��j{|ɴ�˳p.x�G�����9~��"KvO���;| -���]`o*��;X5�KR�m�Az�?fu�o�Q�N_�<5 ]v���ep�ҩ��>	�`/��X�Ɯ�\�4�}�"n��1����r)P!gv��)��J�$�G���u|�t�v�XM�-�'Ճ���7���t$����n�qp���1Ǚ����oZn�q��so�p��1�����`��+
�,m��Ε�AT���p��LGK�}č�������c��6o�\5;�d)���a��Q�ج.�-��G� �j��/~��lm*�hUP����)
������:��A& (��qe}�$�|Ƽ�x������&�/t� ���d�)'�Ak�G'�)t��!���'u�G������K|}��L�>&��68��	%},+��צ��aN<���4��
��V�U�����ὥ���r��l�k��k��9`֗�H��/����/J��_[_�/n��(@	�_T�N,t�� ��ݦr�r$f�F�{����-k�y��>ԩ�EG��l|N�v[��9�V�F���sFZ��tT�Ϣ���֗��;�۩	�>o�"��q��e��2�v�gӜb�䒒��JCU+.�#��T6<�e}��2��� 8����V���^z:]F�gK��(����{v��ၻNIWt�D� ��G�.
���]����CQ���_mݕ��ťMlu9�e�M�j����`G>��.�º���� �L"qgi|9�UH�^ӧ%��`G�Q��.�v�����\���x����񾝮�D}l'����K�0��#���GFH̷��㻦<��~)sݰA��������s��5X����a��Y���(�>�b��Ƀ�&S]�*gz�7w��;!����N�ړ^��!���c`���ͨ�Ee 8C����5����W��Fu��bz��E�OmQ�;*0���L���h7��i1a:qfN|������*�jA'��{��O�rڶ��]��C�a���i���WK���-�$/���V���q�Tm�hY��xp�����w�uzd�~�׿���7�(^����s���$��n���}3͖K=~��0��7��3���^��cuV�B�U���p!ַR���뜓��FΌB�M�����\�Mf���t6<��'4�j�5'v�6��������%�6���~]a&�<��n˵y�KpT~a?��*h�J�XQGrz詧�3�Z�`�{��`Bt�a�Iso�'�O�m�y�B7g������`(�|��B(��p9�l���z�#N�a�.��#��Y��%L��A��O����]ݏ\^�E�w~���(l��K�$�N�G��Sp!��g�H����Q�t$ĽKH�%F�m�X��]�XvF�7C<
�N2�x��ۑ�߈D�*m�IQ���
�d$'�� *�Ƀ����������v�]�4r�d��Gi1�8r��Q�Qmy��K��[2%S��`v�.m3�����ڗ�^�q��@���4�m�o���kT��lq��O�,f�K�iPӷ���,����B��ёe��.Ό�&���1�"w����`DIB�vQgd�碿���)Cj�����U����|���������7d��b �� �'I�>)l
c)���⑯�]13�n�0�z9bjE%��§����Q�!�+�q9o.��~v�UW��a�E�7�kĭ�-���Z�^Y�w��o0bp�Ќ
�.k��~a�S��bd�ۢ1���|��\/����z�Mij���Q����^g����}��u�F��@{��?Od��x�Q<������b�={��_�9�3�rD`����q�~JWˁ��t��9�
�����H5]!�ѓњ��ƍ���Ua�?��,���'cǫ��ʅ��^�>&7���!�CIz
L�K�9��>T�'�.\���c}��mX�<�J@��-ӛ���'���2d�*��(b��Xk �,o���4J�h�)��/K�7+�S�#�����I��*����5Ke;$N�Ѳ�Ln���&YU���J�q���~1b������CT��k:��Zo�4�hƏ�@��|�P��.���nD4��zlK��S+�!p���-���s}��s���͒vȊ����L��ƹ{4���~XT�/5����
�Ք��>}k�*��I��U���(��ކ�Q��p|�8��J���Oi���|��"�$�O	��!�K�eK24\h����b�����AV�n,� %�xs�}�(�!j1��:a�3ݷ�M�>T\`]���ohtl���	��J�: ��2�uq߿2�o��4�\n,�
T�ڵ����B"bm��#��\��ik���+$δy���Ǵ��̋�h.5��2���ތ]�m�G%��*�PW�Y������=�i�A�P�2��ӊ
Z�!��d�`ý�H!������==)Zx�IZ��u'�U�9����n���V�ηmk�{���5�����u�?'�ʽ�-�����̿��M�_�S�X�?���U�`�th݊�x�qW*O@��/qo����^�Q\�)%����m/���׈�U9/���5@�����Nm�*�:֙��I�)홒#-��;���@������K���s��}t?�)��mT%�{oD"QI|ek���U��{�)ϕ59�)�W/B��=.f�����������v��ȡ5�)��g,���PC7�S�S�ap��ñ6�iUs�4}�����<���3!�@��p@�_L�4=�

MD[�P���?�F�2n�J/���V���d�y�_���gy��FH"�n���){x9���3c\I�}�0N��G%�;D�����n�ߚ��x�&׭���˩��yzR��n�gh��|{��+�^)��60�%|�A5��Y�j��=��(��D�A�S7���#,��b�' WK+IPӓ�N� 7/���0��lZ���F6�GP �#�O�������P�?vxTDK�O�A�l���8�꽵}7�s�~X��Y|�)s<`� ����M�?��[���󀽳W'1�Xqv׏�#�t�nY�4�=>�Pq��s�dghpp�d3u�1�xa���t(Z�[=�HU;[y�ɯ	����oȮ\�d�~�ll��&6Sd(&�^�{���WO�����H9��d�/D,�V�B~���v������(zZc����_�OK�����ґ��^zR����0U��7C��=��C&ۏ�����z&x�%N:�g�Ro7S�����L�5��1�!!�f����K>ͫ.�G�ɓm�����[��h]����5�X��2����_��zeK*�������D�hY�TQ�z"UR�M(,U�����1eO-�X���B�~/V�u3�w�
`M�	co��	*�39ʷ�$�,��z{:�L��[
`I�������=ݹ�y}&y',����I^p���^%��V5���B��@�׿�H�,~J�"��>>�4u�VJ�]�kʈ8���c�Yv'�{���S^w�L���v���ʣ�W�.�<�����D]'Sf�a�A��-�=�dЪ�l����f�L��t���Z<�_�m�����S5L,$��J�^��:�#j�l�_-�"�p���i�Rݪ�0�]=ٺӮ޶-�~W��2���iC�i/�Ș�S:"��4z�n�h��˵��'#29���gu�-v�C�7���/V"��O>�un�{fƞ*z��]�5	;O�#�x߉�z�F&K�7��^{���$x�XV��(~��kB̷H��hO���M�j��so�T������T3�?�ĐF���%��뗠�Fy�-#�g��Y�s��/��}�g�ao��|�[�����F���]���NC�ٷT�@�_5���C����(���"|�U�
����A(���r2Oݒy��8���o����㶿t]�2@1��<o�x�O[�
</]l�|��W~X�W�֞� �q���@ˢ��N$J�~�m�¨��ѐw���`~���+�6.�D�45|��AT%���c��6����Q��$ ���������=Ok�g"-���j��}n��H�~B�C�L�A���N��ߜ�I5 ���;ۼ�z2f(��e�?l�6�F�$4t�7K�]��颰3N�Fh�u�[B�$/[9�p� ���5Y���~�K7jF}����+����O�Ԩ�dH��MɌ��I�p~���,dt��dK�u�p}o�5�~�)�sKT��bfE�[�2Yx���f���Q\��Uo��]���w>��VUVi�À��>�-y����v8���v:��5N�"V�}�������O4�%�b��߯�y��u���ʊ8ಁ��e.g�_���XQ��=�z�@���=F�ݳ�k@c�S���6��Zb��xB��X_A%��Mu�qO�ָ�}.E�
���B�G��'8'!zMs2..V`RH
dǿE/P�Q���O�D��n������Tw?!�Ӊ�lK1sl���o������7≮8�u��$�&w�����xv�u�Q�ե_����V1���a��. %yP{;������q�&̓qK����ޣ�S.ʿ1����U�\��h�Ӄ��B$Dބ�m���+��KX�:��r�H��/|\�#��9����1��_�/\�1�xU��	���9�Y$�dM��rm�ȟmabg���q��U��D��e��a(�V`³B�/�8�ک��p�}?y�y�l�R��|tSf���%�cV��y�����u$~�:ݠ^���N�EŌ{��E?U�*�dq�l��8f�=]{Ӕ��'�g��j�:Vs�43��q�ժ��w��-�=Pn�i6����$��$�5%E�H��n���t�'�JPTS���y�	��U��e���=��x=!�*�L�z�}(ɓ/d���� �^q���Q*z�ۡv!��I.SV]}r|fÍ��]��~�%#�SF�f y���z1�A�!`mi�H?:1<es��}�>1��^ΕJ;���Y�������q�4��o��w��!��R��M9*��j\%��.�b�����r�ڦ׭*<�4냡�n��=ڧ m�t��Ω�\?]Ɲ���&{HW����l�b���dr���%���јqB�ʄ�}���ۄBo�:�zOI��I��V�U�.��w���{��(7=L{�^�F]��A����*�2�"����y��ƌ/o[|��H7\�0���O�\wF���-���)y��r�qq��:���)/-�����O,�?��2��ٜ�`	}��� �'����+��5�Nh�gdQ����ﴀ{<��o-���w�s��Wo��P�w6���;�\�q���h����y�ߏ�tҦc�(!q�v#g[��_V|k�N���ٺ�p�f�¾����e�z�>֮���%�P�93�0��d,YX�S?
{���r��H�h
�g�Ohn�Ҷ��5�09i=����r�H6���N�*)�ɋF���}^&�3z�ޭ���7=(I�7�Q��ݐ�[.�8k�Y�@�"Ԗ4��ө���gu��f�wz�X��A���Y�۳:6pxsW&������l3��E�YE��uk��ݵ��;�8Ŋ�w	Zܭ(���R�!P\Jq)��;��U�N֚���]{yM�mp��>y v}oY���7!�ۀ*vW�
Lќ5_�i3���%GA&M�-,Mɼ�Ni�'~�^q=с9kkA{H#�6J�ڍo5�Ԡ��eg��>�R�g�@;aDU߿G�����g]��T"�j0��������]Da`.�/U�[��IB�v�O�C<����0���X�Ge����c�9��ǚh�6ΙA��>]lu_;����\����L� x�z�
萓�%_�s�@�32u��훡{��ڷ��J���U����81�_�\��&Ls�!F�7����Ziy7�/7g��z>x�g.�`��	:W�"B�\��o�=k�9�5�.��q���t6'�3��*v�l��5����Fi��v�)8�e��{��>��87��Z���/��|E��$M�$r�8dI׬Zԡi&I��<����,̄��d���f~	��Gz�ʠE'Ȱ���V��A�1��2�]�Ie�^	���k��z������,q$�H�7~�lt�|���d3r�6��v?d��6����ɩϋ�D0�C9��ߋ�xHe��uzO��4��Y�/ ���E�M�iX��_�za~�zY'�I�e�!il��$���S�Dl�+��CU^Oa]=���>f��Xl�O���}�W�[�ʶ|�6@vҺ�0��������f�B��w�Bg$���,�Fi��**q����O����y�����Ɖ��lq	3��_���:]>WX��rAX<7�}�Q�G�s��f嬹Q"G��Y�3��fOoa�=�!�]�1�J>�{ޖM��c�N
�a��Ԙ�����u��p��|��Eۨ�h9K�l���ή�l��9?{������Y��T���z�6��"i�1Ԓv�=�2m��Y���q~��)��
�x��jd����/X��pBeE��~���D�ܺhg�>H�"�g�,��O��YZ�1iu�f9|�ʙ_.������;��G΂�+:���iJ=�YiM�7	�F��۬Z*�MX�u1?��)@C�M����8�ao�<�r�w�c[:��W1��u��%%�#�3��,�T�gK�*�����e؊p�
��Hg�ZWc�'�wz<�&�n�+�x+P{[8 �
z�=\':�˧:�&�;d�$"���f�BH=.�;Rq�� �m◻m�ZHR�=A 
j��tw�p�VI��՟̏ؠ�����?w�7U�	���A��Du?in��RqT"�ʱ�Bk�
!`�";��L����#?�����܅���7�'�ާA~G17���͢���8Q�@_���7���]:�8J��O]���k�nr3
�Or�W�)���`�B�j���5�P�I��:iޕ_y�����-�qo���O��X����1��J,�gO�-�Z�~-��Qb���c�:�j�e�����O(K�Ϛb�=z.D��G3��<����Z2�٫Z��(���)��� q��y�����O���B�J�d��2"����\r�(��X���%�&��u���)�����:�w�c��y��f7�ɋQ�9�9��n�}�B /E�e�:O��Zͯ��d��%Y1G�~X��ϵ8�8�O[@V��ߦ���Zu����~g�VF�k���u!�0�`2��F
Nc�А�⌑��&lʆ��
A�⤑�D	d��\�mȗ
¢�l|nCդ�'�i��o@ˆ��Ia�ن�|E���A����<3��A�!+P{Ǜ̬wc���@,���� 2����o�at< �>;�l"fxIlGR���H2(ۏ��~�6�Δ��t��h�D�N�^�z`����d��@\apc=�wѥ�:����������L��I�=Af�8gi��ϩڕ�Y*�Nvͻ&7!
�����'�s��Q���dx+@�_�P����z�J2�J�Ω�iMێ��Pu'���W�g����d��i��G'��|9h�q���)����~�T�����`o����@k�c��&dd1��M���<Wp��~fm�!��A��Տ)yy���V	�,��v��aIA�z_@[T�Ts��=.s�(�%3��Î'Lq{�8*�"�z2���+���[�o�4�����ۂǇ
����Әy/��!��ۙ�8�v��CQ0�v�5�W���Ũ�p�>C�Jy���<��/u��ɱ/�ʧq��)S���s����lJ��#�[+�ס�!c:F��[���|�U=�m}@���Z�g5�?�zҕ$F\���T�B��\)Ӓr@�2X�9i,��$KS����^�.�f"�r"ʴ�k��`"_#5g���H�C��y�|�H�҆Þl����/*�؃�Oc��oT��
�A�5�-wy�^=�W�K>�ߋ�|�m��^�� �O��Lc�'��1+Xsq^�I��*��$5��)^SA_���@x�ܠ$ӭ�BR�m/���XF���}>���U���\���C�G�������5�N�ug�>���
t�Xm$F|P}K-
m*B��^9���K(�D\�
e�[��(�?;�[G����X�Rw4`�5DJ��L�+�"����Z*V8��1$�ġgSB�q��0(�3�ƅڟ�M{5{�n���|��������}Fe/���Z�[��A�G�;;�����7�3�a+�RCO����ga�ͧ�[zja���� ��� �GТ�c�m0b�C��І��̍���o	�W+U"���8��T��j���@h*��ZI�s�@u�|K�kE�"~�Ø���l��{��1�ϒN������
3�Z���>��|���9���tEH4ȃ}E�c�]E���k}�%��W-�����M�ݫT@�k�L��EBq�I��5\#j�tY,�X�v%�� ���m�N���0��m١G���+�����r#K�guջ[¶]��`����Eu�5�I�ۢ�4��Dc�bb4Q�`Z����J;�8P�غ�n��0��^`8C�?�p���obZ�u�HY�]]���I���T|�]q���!n�� �G�XS��V�E�˫�U1�B�R[��N��+�z,��Цy�B�t\6@�_eD��,7(��#�Ԩ�;��R����ܴDi[���v�h���K@��)�p�[��ai
!n⛁֯L���b�^�Be��ހ�f�p�}�p�l@)u�!=���Vl8e_�C���m,qi��3����k��{������Hz�O^�z>Zr��4�.Ԟ#�s{Y� k�tf�?Lb�l��9��5�ACV�&s������W;��k�[E���G\�N�Uy�!-��F�M�d��*TyɜA��(BY�)旵��Z����g�Dk��zyul�w(x���k�5����p_����Ѣ5:jĴ&��c}r�d���y��-�$�Ϫ9���n޽�S^�9]��7���3�h��H�,v<�bY��h��n�-�,$�*!
�C	 ��`;�/eO�wVO�[�J����Al�x����+Ֆ�P��|�����'޳V�N�7�����x	��hb5Q�8��N&�=F�#)-��^�wW��$��My��d�,d��Rg������R�L!sW9�v��ػ��~&��X<J͊��b���zU�ʪ�a��{���-_�{�a|Hr�˄(�et<����"2HGL��tSj����7 %Q��:��<�n���|b�7��׮D���ns0�c(��Kp�S���C��ޟ����*�%F��)��
���vB�y���
�̯N����.�IE�&�%����Һ�~�;��Q	c-����t��Öw�}��d��-M�{��n��Z�Q�D����J�i�\GG͐{��n|�F��&�� ߴ���x�r��D��
��ѕ�ٗ�?��!6��a㢓�j�S8Qn��䴜��ю 7��Η���^m�~��j�cr)H`��8_�l~��_���`��&�D7<�~����3��"7��͹hxs������$���Ѝq��t?��&�>>�7i9,�=7��ҕ���gx�!�����&],t,=��Lr����Ex��1b�� ?��zV9�	혞��f*�9^�L=�뽁��J�8!c�d<g��8�ٷ��mܚ�U��Rz;=�G��!�&�=���}a�:Xw���Ǯ��~���s8��&���U(%��|�ɯ�?'%ƽ�B�#6�t�hy����D'�I:�7a���MH�����k�#�r ���짌�IT���wW��>{B�X����I./�"Qո�$jP���k渠^�	����c���9'K�N[nاq�?�i6t�w~��� �K̄�d�]��6��Uw<|��!�o%f���^=��u��a17|� ��@�$��RD������8�n,np]p����p��	�np'Y��*���S$�p���Տx�s��,�u�!��A:��{3=�B7m�L�=L@9�/��\0�r�B�C/��s)��/�>C��|��}��+���K�#o}��V��Iw��ϟ×EE�ڞ���7�LF?&�	hKEv�O��|��󟟁�O��{	6����b��^*�� ���l�KK�4���5�N������A�����w	��_���08���˜(�O�H�aa;p�ٜ�����z�|M�د��!&�$U�bn��e��aD�����
'�-/��\��u�ӈ���zy��4��)�¾%u�ˋ��0���U��#�+h+2�����2c?(��w�.���x;��~�:б�ִ[e�$�Mi@IP�R�bT���%��\�L�F�VJ��]p%F��N�[H��3&��+R��������t����e/0�Hhn.��&?(��������F��j�.�EH��L��њ�b�R<&Q.�)��۝�ݣ��%�%��A�V��h�2H�����T�B�Cg�%��!��*�*�0��$5?���専�zWqJ#�F�ɾ��P��F�һ�\;o5��r�{Y����r]��F�Q�DC{���W���#P��YR���ŧ��.���1�[��0���IѠNo{�li��代�+�X�����J�3�{11��N4��Ę�������K�V_?�>N��Ʈ~N��w9l4��N��t�|�v����@*�7���.�n�f$���O�E^~Bq�� �1��kO����(�f�o�=����l�m�	�#֑	��1�.��|�S����p�6V��n��f������D�Q���R������^�E������wr�ڛ�G�"�y5�;���.��~���뿮_w�>y���$-.BNƝ?@li���ndm@�Ǭ,�ӚI��3oh�w�J�N�N����k�ihܑw�2���m%��b�Y���YuW%�4�ݱ��b�z�u�������|�ud/~l#7 ���Gtώ�Z:��x�C�`A�;h��GE��ֱ8�L��鮈:���V�f]�m���qi��.K������c��=lA�M�U�9�!縯ne�zw%y4�z裣��m���
�܊�L����"W��E����Q	_�w���ѝY���)����MJEr���������yp��7E��G1ji�v<�t*��؊vrdG֏�ߏ2���$�!H5X�VC���؋:#8�͘��XF�n���xKa��n\�0�'ip��xbJ��j��a~�4�2���V�w���IKދ��b+i�?|,��P��;Xڊ|����Oj@��W�[nq��R�
�E5/I���)mX�1훻Go�oY*Xx�}�����^�I�g�C�?o\���C�o�¨(������[�|)��[��$���F?rל�d�=�c�e�D.�U�����`E� ���к�jmpdN����G�͇O+�����3ZEGC���~b�	ryW��J&*1Q�;!U���������#�o=ڬ0�UA���-������:�b�3!!�����m�����<�ӡMB��WQ�Gz��O ��5a^��ʒf����H�*\_�J囻!m�z8s�2�S~��{��"�[���@��=Wu/��UY��;�Z�'�����J���;Р&G�ɿ���k"tC�,��x�H\�tYRPj�~� �j"u��V�W�``�U�^tf}<�O����i��4^��E�'hP"�K���6oiμ�Ԛ�-ħC�KXJ��%E�7��s�n�p�0Jb�*]���b�1|ݩ>�)S��+�o�pX������9��ԟ�/���Vs�Lyu�C��'�d�wyJ�ňTW�4��~8ܿ�-�-xl8ڂ�'P��Ȁ|r���]K���6��'���_s���K��gl�
�w�}���62d>��@�Q���/���U#�~X��["��.CN1�H
��q�V��P�X�p�:��]��G��</5Jx��C�=F+X@�;)�
���O�T���J�_�j�K��50���(Nװ8�������,o�tY0H��7�LK֎p�{H3}�Xu1l�Jfø��|1x��V�����
�⭧u����/>TxG^��,#j�`��|���H���)c�`�+h�W�WR:J@Q������rT�)��yR���CA��Fxr`�����xJF���"��D�[�B�\���;A��Y�i�e(��TX��݃^ 1͍e�}n��¶!�N"��D|KZ-.�;���wd���`/Qݮ5X�yk"�MDdTh��y��	S&*g퇮?:�%�|8{��;���S�@�FdK���7�w^�~���L�?r��*�P���v��7	b��%���Rfz� �� �~�0ӕ���{�^�~���ߖ��v?�y�7��"��������]�P�q�mh�XLn���1;��ڼ���v���-LD���m�����?�iFGb���>�R�	r�t�j�&4w�W��6��Pک�K�#���vSw_�
9�t��*��3�%[���e�ĭ��e�I�uL�e�z;�#~�]��=��|B���w�6�e�Q,���d���rE�G���ЮD�	�F�z7��x#��À�k?�����S������C1?}[�.Sy~�S�cH�q�۾�u!L�O�N�:	�d$�L
�W�z�F�Hb&�KJ��������uGݕ����l�/�m~v\z����N��fr9Z�6��ϯ��a��ɰ����p��k�R����4y�ɷ�ԐlY�Oѧ|Ϳ�������L^iC�,��pF�B�Grl�`��ىQ�s���qs����2�P�K�[�<��ϥK�]�T#�/��4���sL�{�Dp�mQQ�g-j�����]3^�z��À���G���ءksa�e=�>6�5o�H`�Yw,�"BF��о�3g��s��Qb������Fh�̋p:���$��2�ncܘ��g��8�'��h�%ȇT����)6͚C�T��`bQ�<�Hm10R� )�.!4+�&����~���޻��<�R��Y��TP�r�=�).:20����>��}���bʻ��t�@d�簬E�����UW�(�\o�����sQnT)az��O�_M�kL��RjR��� �:+��X�^I�\s��eAҮoׇ�yOw��������2�~��<����S\C��,��r��yCC����:[}�	��Q�k/�2�UN�U�`M�_)��I�"�������(���=��\���,����������'�㯶�Ǯ�#��}�:��9M�RXُ���g�S�3�YӴQx�q�I�Es�p��q�;�����E�Y�z
�OLk1o	=;`�H���K�N[���P���D�P�/��sh�/\�Xpvk7oucr��}�������\
O۫�}�v��4+f;��@ֹ�ZZ���Z)^OwX�$������t`I��L�wFn��.���=��u�5.��8C�8V�[x8�2��8Z���i� ���Ԥ�%>�����0?i��[�<&�n|����;��{tm�>\�.��"p�NtS>��\�J�������د���r@")H�B�_��mN۝�����+�mn�ŶO�K��u�ݫ��Q�ˉ��1]�0t(�˱�Y��txq{~����� c�ǖ�s��VdnHAk��)ݡ���Z��BbG�	׷��q�a^��E`c���QN��R����Z$ݣ��.�j�_w�,B��J\ZD�d߲��&&3x1�Yr���];��u��C�͸����k�w,�	i���w���G�e�c�fnB�I�5ο��m�	�A�)�)��pN�[�
��*[IҀ�#V�J���p�����KQ��ӗ�J�*����(��Nz��](���P�'O��+E��Uatd�2P�
E�8'Hg���hƆf��j�w_������%+�
l!;!$���Z�-r�@�Y���;�h/N"�`KKc����82��KY��T$Aݷ+�v?,��$d����eUK��k����Fe~�{ݶ� ܂m���d��d��Z�9�*�ߩ�x�y
�S����*T�����9\�A|��XY_gY��F3���^��P��d��	9���zg�`��"�d*�όNѯǱ�\�l {�|�ʊ̲f��+jb`{���,�Ԝ'�ЃZ�����������u�
���Z�IdдB�RX�?(r0���"�'�r�4U9���U�9��N4�g>�f�̎T��eD|����,"@il8�!���O��}� U�8\�,L���i�Z�\r�R�c�2�Ϫ�ͷÀ���gR��%���Q�F�Ĥ��B����^�2sl�0��hf��P���ͭwQ��}�!/W�A���a*)���*���AB߲��#с\DȨ�M����������������K;ʿ���*T*��$��v���Ԭ�Z�BFY��b!��o��?�X����˞/e�����h>��:��}U+0~�
�nf�d	���{�E�:�N����U�wxa�,)~��{�P���t��9Y��e�N�힯�nݴc<����M ��'֢>3j3�X�k���e�&q|���(R�o�N��:�d~���|��W��RXa�J0��y��xq��߯����. �T����{�T�������w�w�j��%�}��4t�v�rJ+z�ܩ~�nn?qP?�I��Wp>�#<��\ϝ��z�Z�g�A���NI� צ^ �T}�&qJ����5�7z��8��GY3��&BZ�$�1!�N�q�o��yx�h�&�!;�_�0��9�$�� _�>Y��x?��#ǩm���V�e)A�V%h��g�� �]��,xT�l�T+q_�i2�QJc��c�jx~A���f�x���޿�_�^UC¼����kC�┽XǑJ)�&G��97��n�x��,��k�Tӓk�� �&u
5�A����09C-��ӻ%(�4g�Җ���|��<Gw�k�Ȯ%�j�^�Õu�Q�31�Z,/�t�7JR�)�����6D"KGF��,K����C+�=�6?X���>�i�t����L�0B�0
LG�Eh+|�3�џ�5���T�ډ�����9{�W�9B���Į鄘Ъ֎Ulbd��neY�&'v|�2�o�bL2�y�K���#NV([~y@~�H�WD#�);�픘�������(mZ�BO��R���j��[1��5�BI�_�ܱ�ACg"�{r�&�c�V�{嗃;�
�$��xSjJ���$�J���ڗm�����m��;n��T�Ҕ�GG���G'kF���ի�&����\2zI��m�1b�^�i2��"!�z�G����WCX���8�f�20�u���V����dC�^�kYx�?���$�b�(�"'�k++�(nΒm1PT��hG�W�i��yy�I��,���SH/c���FZg��>>rzQw�B��	�\�x�<7~���됎�H)��������}>�*���39�b���B�6�7l#�v�Կ��q�.oCCV�a�9�dK���L��63�J��u�`�N��E^��_�nM�ntT�c�'���3�a�k�l�0���}8� -ɹu�-ߙd�"ɹ�R�=��,�����=��2�[�&�z�b;�l�5c4�b6hFX���4�M���&U(�t�4�������9w&��ȫP�w�v�L�{����w�2��������i�̀ g�ۚd4�H�1"�`/�  �So�%��G�l�ǻz�m����#s>��:�O8+�a8T�~(�oh�͵&M؉,��2}L�U�^S�:�&�`Vakl[|�P=[J���%���d2�)�?��c�:�L�q_�"�h X�����΢�q;���r��&���c�ֲ�	Btl�x� �8TK6w��ncVR��Q��c<��`L��~�h�4[Q2s��ym䏻	�::��^�l�#��� \x��Y<k@E��՞F��*�	I��F-Q(�T�03��8KJ`��A�Cu���v�l<,���ɩ�jY�km��^�����V<kZ�$�Z�#���e� %�,�$OT�B���L��Di$�s! ��ʹ
���FV��-�)���0-l`bu��_	8$�%�;�S�C�ɶ�ٸ�����C��iΡ>�,���
鶱9
3V�d�٢�!^b�/�b�6_��BK�e#x�b��	P\�|�'��{�x1�ruWgΟ
X�Q';�X�6z�\�:5�&|�?}����n%{���I�Ofc(zz���ي�h�t�n��3� ��\<룇�_�OD=�MJ��qT�t� ����~����<?I X�L[�b#�yN���b�#g��Ɵ�rz0���!B�r��{�b "9�H5k��(�]���{N8�E֖
�g��p��۷�����j8�{z�!5��G��0^y��cs���J��cM���d������!6�%h�+\`���Q��W�AeA܌߱^�ٺDׄc�E���X�'��7\z��4S�m�/l��0b;z�	���xV�ٵ�9E��:o�z/���%�*@x��oS��.FNH���^��ky�B��I�\� �EȤ��b�9Y2(@{2ǟ��9��[9�
�I/�HSm4�v���L+eỼa©��U��X��{{p�Ȼ]��v�9
���#B����Z�9�u�{�?e՚�����:�h�2_�_�Ǫ0�s�KX_܊p�a�Z��j����ߡxP�i�v�;�"�������Q#�salT�~5X9{�D�̱�7m^�A":%���j 3�Gey�}Ԛ��O���$> <?�d�R���K�;O�1�q撕��S�X�m(�sE��P��sg�J�n�=�l��O�|�TzD�a@[{��!�D,��Z��W\��(�1�T8a��c�G(�W��T�'�~	�!���>��?�0��7�)�s~���6��Ʒ����ِǆN�q)�2�����Sb�}�b>�n��4�
�'8pV�=Y��m��I��du����X��۹L.�,v0ϫC��-%y!R~(�d&w&�N����֕�[xJ��ΔU�F0S�8�RZ��d�&qr����z��:�^��F�����0��0���,vq��� ��a������^��Y��B�0��m�^��k2c�����F�H�))c�(���(�����T���졆BTY�����į?�XT�1����ؤ�=�.���+KN7�y�C���@�.=���B*z�h#gϸ�T�Ӕ~1�I��&�3E�)`��FFy�bd��S�
�@�"�"&f�H1ʗ�@��61�\��/8������r��c�����^F!NJ�{�~.I����f��s ����|۰�����^�W��&{��L�U��/(r��=e@m�?@�(�:��D&�݋Ђr�qi�u��jY����c���htm�<��B�R�����<����z$bL�P���|)��e!�S���0d5K%X*��Z�҆�s�jΏ%�)_�Ig����
�|T��WD�FuĒ����%�0�wR��3\=��I�)��Wt5,m�^��n���s7�?a	�T}7^��0��D����wsd�eN�"pe��W����ٚR�w���?{~���a<t��
�&�w����h���V,�ش;�Z��<���7j��p�Tug���˃H̄��0A�2m�0bH]Q�㍖�Tu�a����<�ſ�."=7r!�`��w?�0��~j�`��������sv�®��N�6���'���Qb*�R6F��H�?�j�5����I׬;�G3�J%�G�_^@��6)[�:&+���-p�i�À�m��=bs�{:��]�I#`��� �Q�+��#g����"4f���/?iO��_�$��~�����*�˸1��?D����+Z����Xb#\����Ё��#��9M.�C��T'�
tC���">�S�U�M�.Y�n���rY��1�IǏ�=c)���\Q��te�;�U��4T���O�pB	�H������/o�����$�Kq����ʟ���_��i2Iˣ����@U&��)���'��QO9�w��g1�\��'����%Yp�Ȕ�~&3?�K�uE���Z�����LK�1�Ӯt����'Hy�d���̎�� �줎��Y�a�����U|�����	B�!I���N�����/7~Lx-k�����F0T>>��O4��, ��n�0kY��o�arR�7|������ˁ�x�=9�3�Nv��תe��P63�t��bD���U��L�E����M�#)a��/_��.%b-��ɡ ܽ�%�t�$~4�>~�zx)J8���1�*K�b��xF�BΆ���g�	w��t�� o�����݆���]�6����e�aGn�uh�яٱ��"���`0T�}(-�P���i��ݨ�����]�v���.�>�p��p��J�D�Rd鄼��2�ԋ�	Z�y��0�>/W�˔o��]0�x�ozc��	1$� ӏS!?/ig�4D���Hs�y�Hë25��6���T|�_�	.���T	�n��|��+�_��rb)��ko���E����/K{��-�sH�с�n��FY�Y�-8~��W�y��-Fȃ�9�Z�+��y�Ć��F��dSu<�	�F�&��F�8N�tM�XD��YV�yS$��-��ȿ�¢�7a�����J�a��s�Z��)&�HIx�6�	�;��z~AL��R��;��`�j�}0��\%d��`���q}�y��pٕ ��Ǉ�5p�#��.�}���^�&' ��R^�L�hW��I����t��l����
��ҋ'��sX踞��C�0�����ZkC�F�;�(آ�'�4��[q�B]��ؒ���u"悼8Ki������BH��z(�_�����mш>
��>
"�O�<�Zx���ڈ5�VNvVp�j���k�����=g�U�VV�1 �,l<��2yG��2r�E�B�8�X����lb��x��m����r��-�W�c@��}9��K�UJ�܏�v;k�'v�Fù��|1�Յ7օ1).�|ٲ0�9�9|�J���2�;����o~�
W2 j�4��?�}I[S���F	9;���Idi��.0��f�����CF6F�(��k<U_��B��bŚ���ݺ �}��~ e�T92d��6�h_HR���`a�~���^�c"�Q��(ah��T�w��U����d�r0Sb���o�� ��j)��$=W���a��#|l5��͈����3Fi�11ߙ;��I��ُy���x�Uu�ηͬ�����$C0�����,�~�ʀ!w.���رTyjf�`;J�"�U*k��m�a�#��K��'XK�Z)���Öf5�8�8}���ߋ��������$�`�����K�c�5�����џ��:�Z�x�&'�"�	(�����q���G��:pEd��I6����R&ȟ��en��ޚrxb��J�N=�kѸc��3RH�
[$���,��93J�ءUq��ĝ)O�0���`
y�5�R�����;p�-�$f�TF�V��p�4�Ʌ,txAa>4���T�Q�H_ �6@����ԑoH����rO�!?�ƥ�y�?��A���g��V
���� �L��,זx���-�i"F��;�*��x�@����F83��?�(�\�J_jo�M
Mm�6I]A1��̲��;hA��X~=�ƱTs�F׏r��|��o�o��gl��vV!0�;[6{�!"`nE��7��X
�[����k�*p����#K�Q��{8gi���ap�!�̾�V�Q$4�-�11$�0Ds{��r��'�܊꜠�&�ؽ��C�:��%�˻�?�����>�{W��d�-'F���d�\_�4��������r$����;���p6�}�b�i�15��%ɩ��F*s���7J�������-݋��ƌ-���z��Ȣ
����,֏Z��b]`���8 j�NJS��l0�����5�1ޔ(r
�!�;_��pc��9w(�#�}�Kb�E���GA�y��f�� {x����JD�Xs��e���� J"r������m�8�(�6Ȉ�8�i�N�R{~+�9؍[��"4��5����+b���lt֓� ��4�f����=�aaQ]���|��^�]6�:���RXjd���rIT�	�����1��|o|缷(�W4�����&h��k6��U_�k���_׻,�}�$����E�n[�xo��p�V��)�c7V�}�:);�.��qhK���a7������b2��#�!�>Gf�S*|Y"��drJ7�m���ډ��8���w���ܞ��O�wB.�M"��>��'�-{~�sE���Wp��K��0��������`^���"q��2x4��j	���C��$�w�3֓�:{�_��'�N,��5��6��ep���Y�~-CV/q�(th��2J5���2d��:�%�0YJ���c;�Iе���wM3��zxXc����<�N�é�4o�˟�~����8Ԩ4���?�y��m�8�>jeMA�Q�n�w�_q�ֱ깧af]xnCdg�s��ĢChW���DЛ�؟2(�z�$[9���6F�e�2gYl���];#-��b�3�����v(�H��}��PՋWs|�Y����;�����rd@E�I�]���΀��OY��o��ec�������ߖ��\U���w�)�l(´�:L�����<�[a�yI��x=5��$������g�
�ȟ9�'�?��
@��� 5���ɐ��@.�fS�Jmo�"��Ns�\�;��ڔ=P�ao��� ,R�Lpʭ���b�B�j}��A�+���L�T�p)*���R@�H��ߊv��(�}*�L�m�#���L��]p;'�6��A�X�fԄ��_q�{==�
�:@	�_�׃�?E͂�#OL�=��|cEh��˯�$���G[�W�w��Y��'�*��>#��M߈�{�(ߕ ���%
yߕ��j(�b±�Vq���E˅�::YK����׳Xo%�����X>� ů���p�"?i�IY|�b���ǲ��$�/�$��T��~�V 4LG$�����F4�I�;I��uBz+܍�_,���0 ��ͯ��V�� /�4�a�\aļT�Z'%F W����}��u(�)R��5Ʋ�c2=�LT���a	�%������ɁI!ư�̲���v5f�o��nu_��}�d�2Hfm.�MKv4"�뽼R���꾬2�(J���l(���C�G�`<�q��J�z\`%�����=�.������䤪(O����L�d�D9�>_���X�'?�{Y�( �rg�ٮ�ˑB��޻�?W�����	V�;�ݫ:��$﷿�˩�Z�.\�DS9��C���%ʎ*��}w�Q���P�/L��QȢvb6�!x3��o:��|z�Uz�@p ;���;�Q�l,�gi�ثZ�L���޿x�����z��F�a�;8Bw�t��K�F�u�6ƉE'����`�+���F~�Scy�������ga¶�1�I�w��z�I�8`�ol���{�=�)oX���L���
Ÿ�Z�a:.��Hø��Y�Kd���L�9�u�YǠ�v�;�@?����}�}XH}�^ݷy�Չ�G��#�{/%��CV�a����vٿ��
�s(BdK��?RGB�3��Ybu�A�?	!�H=ocYa�����󻮖��-&�o}�M�Z]��)E�EKGr`D�y�NQ�N�5"�U�!��o�F+���"[�ܬ���;�PZ�P�oْb��Fj�}h�~#�3�M-�M8ș�f7������|8��LB�m�U��ɎP0m�޾w�
����ͽ�SrL���,LxΒW5�PX�eCl1�7�rK nHTeAt[���%z1�Rb���aSW�N[�p譪��a�t��Dx�68&5����t�m����GS���8���z �)q��)J�@��4���;P�����qHZ�u�N��,1�\��w]�ab��(�{ ݁�f�3���
)�|$���<k!Y�!6؏U���3J��B��3+Z����b��G�9F���mx��j�4�m�l�ƶ�ضm7�ݨ۶�4�;����u��Yg?���:{�3��2�:I��+6��o�-�gQ�Mߌќ��f֎Zk�m�0OS��[^2��� j���4���o*ҍGDN������zl�����Ȥ|s����V1���3+��YR��[T�j�����w�UvT7A��B����A���?� �]�ښ����H�*p&�5���I�q����_����Z��|8-ʭW^{�h�%{h�D�^�k{�A�D����#��/�a�V51�39JA�'U8����P�9�ҡo�`��'��p���`p��\�4ŀXɈ�>�Z��
e�|��4y��B�SQ�������r��
���I�ќ;���6�����Y�j�$&��xe]�V�pY���5g�N��,�ݘ���qP�y��;>4�����|S��������-���#}�5�5/�[H�J��G�%FF �0"B��S��vթNO�oHKsz5����g�j�V�M��^�Wܛ6��4:=oNX�t��#{�t""�(��&��M��;��[~���8�1��j���	Υ��%b�Y��CCڞ�U�����J�η$-�mL��p����7)�"�z��t�O;�^>���Z2���8�$ʡ�]�Pk��T���k�A��B�.�m�d�??��Q����.�\����!%.y����`sL���#��<�jI���*�����7;G�x������ �$�Q�
��c�c�_�3�k�t��G�@�D��OK��y�����<��1����$��E�;:����X����~X*�Q�9�0`M��/ɿ�swӏ�.�G�Q𱠀(e)�1��Ω0FS;9 �?O��p6Z�W4����6�1�:��U�<O�)�o��O���v,�����QlQ;�d�2[��b |��P��E(eG��@�ƕhVs	T���څ�"���f��m�ʔ6����N�	'e7�ho�MA�:RO{L��LA�_�wj_��0��X�
!�Q��Ρ*ʱ1a��8[Eq�z���z�p{��}L�;�J�尀z�^,
 QY�{!	O��業!@��	�����&T�{�{��{n����Ϡ��H�
rV|-��Q�)���z �0�B�t�׍5^��Uv���ueP�6PeI'V�Q����1i+��>��*,��pZ�7�'���lTP��V� i��ٝ &[|���ۿ�G��z��Oh�]3�H�}7J��.�z����r�A������Ө���oP�=�M�Ik^0o�o_j���U*>&��:��J4��\��Y�0H�m2a��|Q̩��jsA�J��M��v���kd+�6�LJ�{�Z/�P>2-3�.lўSD��בMc(�����-Œ{����$�/�e.B}��S��Ȭ����)o�{���̶��tY��hw��}@�6��wM�kFz�e����#(�5U��S~y��G������%5�wf���i6��!�)R~/�X�M	|m�+�u4����*o��&��|10�{�q�5��Q�1�֘2�,f�'��߿w�CP��%�n�K�ftY�pc�BZ�i[q�c�I�1�'ڌ
�i@�N'VR��Ŋ?\�/�/r ����h��I���@� �=�Dً}6�hY��8��h\�߄�-���	
}_X�'�����x�����o�O��wkw��e�Q./*�x�r�J<*�u�J���P3 ��`��q�mJ�D����)]�4NDM7��G_��oC�����:��(���.Ù�����3�'�"L��M�L�m�1�o/b}YYx-mI\����Τ\`'=�Q�
1ވA���ޚA�ۆ0�v���������aNg�^��0��y{����w_te2�D[�9��}|�J
LU&<`�PqA�ˑ{uq!.:nX�k\3�U���Q�N�đ����3r;l�E��{Ӝ��-� ��5��x���|:��}���T䱘s��b~�Z2���^�>�Ɯ�`�Nr�B��{q��s�B��������b�s>��G�MC
�6��kY�O���T��)-��g}%JR%�����W\�`EYb]'Y��[�A�f04m��*��d���]TxDn)|�����|ǔ!/E�w�'<����O�d��(�uF���b�u2��u̫�q��h�c�����
#���Q7��&�ۓ/�[^^���V��8{��u���U"�S�Y��������Ţ�Tg�̹�(Ć�h��AM�t�C���cW|��;�gO����U^7��k�o)`�5��al�W���F��3����/��=�Z������f
�ל������ƉU��k}�P����q��ks9Զ�a7���OW#>�G�U9b�*L���9Fk��!s�q��`t�+B���nE��%5E���w�-��/s�ݾ|������lbmW�s7����&�	U�^�v��!�G]�]�S2����b�d�;�j��:� �>��/�l�TDV�b�۴B<�7f�+vTY�U�d�ï��i��cѶ���'�)�MY2�B���lm�(EI��Ш��+�l�Sܼ�b�ɚy��d@�D�(�%���Ny	kq���%�a����*}��_��waZh��T����u�ٹ���bo�xJ�F�pyW��L����������a �@RvcL:�K���^�br7�㫸��Q�٩x���nч�iG��lb���֖$�Y�a���)��A��u�F|���� ӑ������uy�Y)*<'�;���@�h\�3�.;�H*��=����rԑj�"D�ؠ�#A�"X	����j�*t���5�1���5L��÷���8V(�"����oz�1�==IQ�����EZz�k��W|�g ���+��wG?>�$tS�C;c���6�`�
DO)VȲ�\��;W&�-g�HC��E`�a�7���m�0,c��X�}�k.��Ґ��?�}�
"���|���|̞��^�ETAhnC�0�5�n.�yұ�_�1�Uh1�.c*�^)����L��TDg����5�R�`|�i&+q�2/��5��J���c����P�	髄QY߉��~���.}J|wSL>�����A:�v/���hw�/�e�-�O�|N�:��`Ir��+[]��v+߭��?ѽ�hE��Tv��pI8E����
I�xFM��^]m�x�51��hf_~�Gp�ء(U4�+R`��ܰv�p?ܛ&&7/ю��$�y:�`C��_;դl�����)|�ii�v�ʤ�qBQ�'/�[����f�`Za�s����0�&a�~^t��f���-}��'}s�RkCӭ��\g� S	���H��-e`B6x�4���Tؗf��wU���^�T.�˻���'�?R�ԔQq�h�U�b�V���su��9HG���!��hQD1p��Wq�K���H�����������C���-�G�xL�����v��g��>�	��mBJψ5��>^�<�m���zg��cRYi�/\�ԭ���[JG^!�6��a��U+�֞$��	��ޱ�V����hȨ�-�L�i?fV!g�s`�oJB�*I�4�b%P		�C���K^E�Ȭo��v"��e�դ<i�8q��chH�~��n�{y���1�~:tN�G�����DhOJ��9���4���o�=��A$�� v%�}VVQo��d`��x���s��v���pwCZn-R)E�2T���>\H�=�3���Z��	~㒀�%xyVq�K'K�P��1A�zd��,�2u��ݢi�Ƣ&vY7g��EiX���1_{�i�`{ik�%�
Ig����gXڔ[�5"\H�]��x��7;�mnU%;O����R�Q�p�!A�Y�k�=4X�Έkæ"�"F���$ھ���O��F�����ߔ0
�|u�
�������W���L�s#�������������5bu_�r��ʙ��3��8<s/	������"����V�0�Ĵ��̹v�к�#5&���`0��be��H�,��i�pٴt}!�YH�ﶃ�
"F���{#�9&�<����奍}������o��R6�xy������t}�JR�!��	�� (t����������l3ΖCh��F0��ƾ[��MK9%��U	��d����#�3-}��>���P�c����f�ӯgf�r�*�U_q�������Tg ��")���д��=vž�*�sIY��C�r�����~��?�P[�v?0;����:�6������">(d�>-�}>ͻ��D�P�˲:&%�4��e|��k��{����f�c�/`c0ΰr����U,�\���:P~ec�@��G��UbV/�_����D:�s�r��n͕�K��*���;�J�4ڔ��y�q��2v���Ef�\�Ƶ�IF|�����U�X ��o��Kl�r.޺|2��ՠ��ˑW�qy&�����%�\�wx�	��]���������Þ��_O��w�I���N���O"�(:�Ԥ+Ӏ���LCt��oǩU![��=��0R�Vֹz�eXF�CR,���I�-����p���b���h�S2��d`#ݙ�����V$Ey�,��9~��$��,��ۏ�ԁM��.m�a�IK5{��9Vs�[��"��:�D�� d�,���7]�W��c]>�6PԜ�:ͧm�A�v�?���[8SH����+��$����G`Dɨ����j�H��.`� ���vAcWI�'�$s���olS���b��rA�oA|)�ި�\�1��f}���'��պ�"�(���?���n����To�� ���H��tY]p��V⨿�N��mIEt<�fֆ��L�V	r�Vꤝ���i־��ݏ1�����%Hb����sy��Ss���ze��Jt����)�|��=o��ݡ���4��`w�ҟ�����D"�ك������х}l��1��p��wd󊱻ܮ�J�q�gʓ��n���Ϗ[N���nR�U3���#�p�ق9`Uˈx.R��m#�~�CEj1�p��6X��Wy��2b����`[K��D�&�eC�&�si|�M����@�z�Y�F�{w)���]�+�:�3�OI�e}��*�hKy��,���#���߅mD��q�CF�É������c����zuc�Kr9kW<v�~M|"J��Dtn��	j���K���J��a�N �:v��yP���b���9F�5*G��X�;ք�Wqt�
B�4W�r��^��NX��p�><b?�0b�Q�|\�6��[�LDV����⊘���e�)"&[K9�H��}�,��������k�2���n��i�����O0zkR���wU*t��J�~y�[��Xc4�^?:�{����3����(Wإ,ZUO�8�G�p��s���W_�XU��'���`�5��Y��_~��S�y��W#��<���4�U3O�J�C��s8^z�蒶
�=V����V_��/�0>U$��]���k{>��!C���A�'H���I�"�(���G�;~�%��˛��a�vlt�|5�µEf�} ~j�@ĝTh�i�m�̂�ko�͈pr�v���vY� Eſ�XmF܇?\9=V]��S�ߦR����>"^;��'l�;�`��1�a��j�B QwKp�w��������,�b������?}�5���1�W�v�(�N/L�%�W&[`���M�y|�h_w_����d�N��-����Ը!��r��n�8�l��2�r�X���$��#D�/%�z:N�r"V�\7	n�@_��F�����&�N� PZ ������L.p/l;��5��X��d�h�J�馂��ǻ`�GϺhp[T����C:���<O��%N��5�������k�W��t\Ŝ���eD�K���s�
;h�������3t߾�&���8{�\������S6�0�3�*�N����H��$�x��AQ��]��XM�[�⃿�v��ʞ��I���B$��2���Q!�ѴOM���''�*�[�����2���x��]�jvd����O��%�¼�:$R?�7}2Z�#e� ���$��S��?����K��w�{7�����ȶ�����F�uT�L���v��Z��~<	�����
^?c�p*��^�u>M`�j�OԢ�pc�E��l+"9���_%*%���+�=�F��Y�(�x&;"G���8���)�to����0S�!�`��0%N- B!�tj�� �/A���8��cVoL:�(��r?s%j��rf�e:��TQ%�"��*zg^F�Â����Z��!���Rtz'UR��f��5ifFR��W�H�V��'�?��Z�mЗ���9��Z��4�#[���ɓ��D���]d�?�
?�]�>y��d?�66W�O��$��^����>�ƀ��+duu���~�B_�/dK�%��g�;-Н���I(��_���dn�
�]���Y�u�>�6�~���6�ـX[�D�5G4�v��tJ�NK)�=�Q�:�N�`|4��O����̴E|R#��ў�)?���5=C��*o�ä�E�gF��c ��	�z�C�g0�"ǰ��6��!�{J������F?̸��}7ۋ�(«����u.��V�~�s�26�/6��7N�
W�15���05.n�����:��`���^�r�>"W�A�
aV��n��LR`ͣwݖ�H8��VH�>�݀j���P���V�C�F�����2�	E"C�U5)�M�f�J����=
R��F�.���Cg�'�%�����m
A��W��/nD�i-C�S�����D�JL"x��q8B�GV1�c�q��3QF\H�Ϯ6���b�RݘQ�p��4j��6(��"���֣��0��OW0A�f`�3��f�ݤ˗@5� ER�˖'[��T2eں�'\�#�Q�48q����������w�6�!��$o�nbT'H��B�C��όL�VeXy��a����RF�iaԼ�N[��$KNd�������}��� xq΍���wG��r��P8go��jWCven&���BC6�0S��w��a��"�$Ү��Ŵ鈶V�a,<-�����7أaf��!���{>�q��,		�]�{���ЕD߳����
+��'�D�/iQ^�Ά~�K��W�a��	��	�X�����r���u����v�-�})C���uh*n�^\��_�sg_
fj�{t�uRa�֓��NU������y��d(��Dv಄��=���ؚ��Vɶ�+�E��r���qq&����޷� e���n��C�*�yK�R�j�Jl�jcL��5�.$&zy�T�4�H�d6��H�2hNV]M޼���٢X@�\����w�C���N9�cB[��w�S���^y�B���wS�,F�'�c@v���w��B�D����U�/mS~j�����ֻ�9C���BDd�թ�oROBB�ٗ�騶ӏ�!��;�f��fN��N�%M�X������̗���D'���J����M�u�����M���8,�|>�`�W��6�t���������B��"��Di�ͷ�1A&����m�.�y���"7�_���k�Ч���y��q�Mה,�D"��4d"���Y�����M�8ٮ�/�M=���z�yຯ��8i}Tx  8Q.��+<�U����n�H��h ������/Jz�! e4�A�t�n���{�l)������l�kCĕ��8OVWԭ�N@�2�*+\��I�/u5����?Ì}���Kh�'<[��7�V�����o8�C/�M����P�����h�����2��;֫����\��a��(��A�3l��*x�
��T=y-���f�ݛ���	�n,�H�_H��WV*�sl��4,N��+�P|�
݉/d�kvYZ�?kعV��ݭ�.u	�x���'L�� �X(0�&�6B�\\a�{���B�_Ra
���./�)��q��� >T߇��6��u�pӑD�8`�� wI3,�0N�hM��EH�MY�rp'�|�ޏ��k��z�m��<�R�LJ=Ӈ���F�\ �������+tێZB���}[��X��]��#����TB%W�	v���%�i�2�7�1�@�=L�.�`����>FA�h�J����s|68n\����R�_%j-�b�]���j���y���S�#q-`t��&��9}|X�OCAtDn�%|�R��s��qoVn-�eމ��K�&��q��Tּ|��� � ڇG���%z�y��6Q�qbHX�.���t���%9h�=jW�m���XlŶ��D�rCre'�e':%�/]F`�����"�)؂t�"�jT���D�� �" �f."��	pAUE{�= �Y���	R�0�J+*�K�4�����V%Bv�{bs�~���!Qc/C.�V8rQB7�9��A���9Nź(Dll��CCILO��E�x��a�2��xi��)lr�,O�BU�����J�iP߂��W�a�@\{� ��߂�/��C6~�BbE3�����k�*�R��sH�WY0�Q�����|G�8	=ȗ����П��佂��u�����������mOg�h��o��O������3W���K�!�-K���0◛"���M]+ h�+9'�jW%g��ua5N�8L�X�N"$���X2�����T��8�7`+��ug'D��?���.�u:�GL�\�qhъ$�U�ΰ�k�ژ��cn�>��hs��S�r�*H:�&$h�t2dX)����.�
�j����W?NAG�&VHL�.Ŵ����	���%�����0t����0�� ^0�7�i����qF��V���׋�;�/���:5��t�wK>	fچ(��} �fB��U�|>�n��bb��%�<��y��6ޢ�[�L��?ZD�qrK㲫�F���$p���)��ѭ��Ѓ!�4�0�љ�w�4�K![բF��X��I���l���"USf/#�8���E{�&f���8�RB�v���7pߞ����^��d�J�9���S�T.�];5�"�j6c�;ߴ6լ
`�^s?�a����:��u~���i��a������	:~S��q�>��*���h����F2�d��lO����oU�B�e�&sH���N�k9�	M�����9' �-���׼/�@�q���oK%o�	p(����!O�xb�z�T_)�2S��u�F1�XHFn�`�Ī��L�kq��``����,(^A��+>'n3��D.t	�0��|�.j�~,5��L���m C>�P�l~�������4ߚ��[-�O���T�?��	B"	h
p!��!�d��'#ئ��hN�ݮ_+����8�[+�r��W)��<M5��\0X{��*p�$d;�N:����6_��ƞ���2	�~6��x�j�:�7�o��^ʰp��s�AJ�kc%_�@ȪjM�\�If�TFm�E�gGV0#��:�ӽ�|#L�.-� ��a����۲:0F9K"�r�Z�l�&�peh>ǚ�K]>�u�(R�nv��Oz����x��D���{�~Y����ϴܤ?���f�.��P&�.�+������n��c;j2Et'�����F \#�i��d��6��cju��6h=}d���G�Ą8�=����ĴؼFj��0�t?���0+��	�he�ʓ��ط�
rd���;'�i;��Q�zb|�vW�݄�� �X�C�V,�"/pg'��ff� }����nv���s})�w�;&!�y���,CI�(��M�@�N��U��H�u�"4,���/S�f��#`�ɠ���nS;����mKi5��{�X���&%�W�}�/�y�n幕�%�)�ώ��'R|Xb��[�����f@�q�U�) GnJ���?�����r�?q�5���Eq
�Co�4�i_%��<�q�Q�Pn��zt��Hq}l�a[å�1�UM����P.[�P2��*Y�'C���Tj!o���i����+n���~��U�&�h7H��ȉ=ԪI�� k�z}�����p&�����y��F�Sqf8V7�K:���쑴��Α�����W��dlbZ���D����z��4��Uy�կܼ5T?=�q�V��mp-U2�Ǩ�����d� E�P?G>pY��f�TxG�3ɴf|�J���G��j`>h�����K�^�(y9"1���?�.2���C:��v��r�S�k��a0 �뎠f�pp�g�՗c��w~q��B��x���]ؤ(O�Q&�.��ʗn5�>�f�!�����;v�o&����|���M�)N�"S�a-#(��: A,^�/�pf����ƪ���,s��_�x22����U��Aq�L�ƃ0|+�v�9W�����DT��]�^��#|X03�G�d�h{���89M/��l�}��*H5�^��^���"�"w�|:O~[ӂ�p}�#U�?�OK��	�}]���z<�yê��$��שq5��W�B�6C�)�W^t�8%�4~ߧd9<4�*�T �����Y�&���wE)|mJ��h:�'�Z�=������^+��v!"�2�N 5�+�&���֚)_~0QA�h�x8�[H(q�!4�c��y �[��G�	��ÙB�M%�6�ׁ_��j<���Qh��h�̾=O3=z�0�����}6�  @]��S��pgڦ��$O�`VW�!4rD"��y�@����`��WW56U�l�EJ 6Ѷ��6���ϛ���*��ae?�\ �S��ϼ(̼8�E�	դ�}�.y���6��kFX�mA��}�r�@P�{d��V����pr���&<_����z/�c�SD�`h�q{���.r-J�z�����������H�WIa��Kl�F��6W�Fg|�U_��-=Pj����N��ul�>K̙_MAI�v��p�����e�v�n#0&cE �5)OK,�b�2~*�%Cg�u���'?���n�jD�Q��U����V���U�t���lG��9+Qo{�(��wW�&�s;7g}Qٽ�Ω#�a��3��x�z��8A���i�c���u���	h�m����¸�S��%q���A��d\c %�W��"	)ߗ�N�}ȕ�����>�6�)0^�@��M&�P�x��f���z�EͭjV��Ɂ��v1��T���|J��X4�x=<
��^�!P@k���}(�yH��7���ݾ��6">�������X{��^�$f�`�sY�:�V��Y��]-�.�x.�jP]��ڡ|_v�]u��)a��*��e+��_��J�%c�և�G�	����a�Gv^e^�jF:������8���ɩ��w��9�ͣ��N����9��b
�w�~���q8�cB�07��G�߳ƽ��GA3FC^���N��X���f-'��v�W� "C�v��s���Ǥ�w�{���
/�����sۼ���_1�O&4(��� ��%jw
:!�����y�7=��y�3I'x�+� �|d�ݿ��
|����t��?u`���qy�0�����mڲR�$E���Hzx�M=��/MV˄E	鑲pV�g3s9M������Kx���F���žQ����X��H���5���`��FĨ�`�,�T?ٛAFR9R
��#5ڔ���P'�v\dS[q����W*��Q!�"|�WS����9�lfp!
�}����7B���u���F�G+�s�^�n1`�Z�߁�ߙ��ԁ{=m��3ŶjT�]L�Hǻ�C�L5�p=|h��ټ���mT�u�G����?�����5���<e����o۽�5p�݀���68Zｌ�쯬�.]���z��G^+�BX�BH/�q�sυEo�HL�`����dr����7�d-�vx°+�M����<�q�)O�r�b	|ξ��ɦZ��'�K�[]FYd8d ��Ǳf
�\!�"[o�$�_2A����C K���=L��x���:�S��MZS>��92T"�0���V~RS��
���
+�YZ��F��Z���=Ș��Re��V��=���Z��9E�L\ţB-�?�I��[�w#/`Dwn��$�>O� v�c�0�jS������6���W��7��20���2��?_���-�O6�f�1�;�rh��V�~h:��O�c�V��`I�6k�А	c�x3<����ąM�Dr�����&���|��/��wM����'�b�H�I�����4ߏa�D���|1/.w����\�3U��
�Z�*p��P�-�r�����h�j�)z�*�;4d9�!kfs�	�&s�6�ͩ��ÃTO�^�������ogZZ�r#6(��]J���Qb'�)�Ut��Ლֻ�����Ir���y�J���~���n>'}
�Z��
�O��c}�t-��Մ�� ���<?�)�F9�o㊴u9�;�K)3;&��⛞^�+uh����՝/{�������B�V�G�M����_��hc�=�\�z�//�q�:J������zA�2%K�6*�$R�q���`a�x�]S=��D3�\*^����	|��c5��=�u1
�V���5����'h�2����:)�����c�<\	`!v#�s����g�V�Ţh=����g�����|j�x[���(w��`c�1'�	�;J��
�5�����Ө1~ϐ��ۧ��-�-@~P=2m#K���n����dY�����:-3S���m��0�o��߽M��hr�o���0�p	������~R}w���<�!��m�v�ċ>��0��p�bu$z!�^)��a0�w��GG�o����]C��z�P~9�\�<��S��o~���k�A�� C�na���a7��UdUV�<Op���xJ�N���v�������~�,�H��&HG�#3� ��}�M�(6|͑��-��?�� �5�dna�Z͐���dT���h���z�d[_�İ,�WA��a���2�f��053��cu��x}Y�=��!�.���oQ;��/�6!��Ul [�"���{��T�։w�O�,U9�N�������)�k�r����F���鋣�2)�U���Y*r@�C�o~�?�I^���u����qM?=��6�Y�VD��z��vCxNꈴ���^����������JF��x(K��cL�i"��&5��2��Ö%5�����a���up��X��E�峇`���p�5P\�~>�G��W�!���}���JEcLLڶmʦ"z?���@W�ON�z[��jFk��"�.ʧ4�Gg�����R�#���������&w����X�v�<��_�V��[�\����=���f<M�r��:B�v���z���-��B�iƕ?#b���5:]-զ˓�2���W�4�ch9�)>�t�<�iU���]���s6��k�4�ϟ<�x}���
k��t %I�A�A�=��xt���4	^��XQv�v�v�L�k�A�x�A��8�;�Z�,#���z��`� CV-���<%�=@y<�l6�V�B���)��_��!Ӎe0���Z�ï�ZEar��'�؋zf �."�|��0d�Wg����,��������//>�JՁ36Cv����>W:���z�b!q<�^��*���jed��H��p�����5�Qs�!B�Tg�PG�a�ː�n쵽4�XYB6D�8��6bɱ� ���ο�ѓT��d��yhY��i\ 7�v�l��������sXƩՕ$�'�������?{�,�����>��Amn�͟p��j&N����I�		!cK@���I��V�3��0�MYa3{������S]���&M;Bm�i����]��U�̓io� b�%Xf����
��*�񬺝sSo>�2Հ�A�rB�PI_͸�.�S�fX��(�a��{���y�y�J����\��e�x������m�$���^�K�<��)6\���������od��ր�ŭ��Q#��W��N��˳~��6��f،@�(Q(���2�y���|�/���9��b,��^�5�3S�,�R+�"�qX��@���Z�����S{/5{��7�=e=щ�<r�r:H�����p7��k��b�dg�W��a���#�n�W}����|�#O_eR����Pb�rmh"e�y������歸6~>VH��7�#���M0�'�g���d�1�K8�ؿ�v!���$��@��H�?6""1�2\��yj�ƼT]Y�Ѧ��t8�1�ߚԵ"ś�Gd^�#�Fp���׫]y75{���9�������\�#�V0�N��։Z��6�T|G��i?f8���t7YV$���
�����r�x i�v@�!��笆�0E��o���׹|��oG�J��m#u�Z�T��}�G*���H��8Ɏ&��^�VMY�scW�`�0��$�3���[�G��A���X?B��&A��s������苸-2#�Cu{1ϩ_@y5��FBa�p�Kl+P��Z��+�E��mau�4�g��@��-��������̆������Z7pW�:v=3�`��� ����=ڤZ޹���i�LtQ���7Gg��U��>Σ�F{���V�7����w�0�#�<ըz2������Ơ�Vcw�˨����)��Щ�I6y%o�o�!�;U�k�bE�-�^U�����}.���|�O������obo}��e/�7�cm�` #�+��ԏo�q�L��]YBJ��۔ld!���1%�y."z.��fg|�+�	7;inP���,���h_�,����G�*��IQzG`���s��"}ye�Eռ�����S�4�=k�%D1+��E��U�f2o:)4_[�����[�L��דX��ڪe���NрHm![9TUǊH�WP@��۰g�x�M�6H_�W4-��u���ˁ�A[���Kq�H�wX
���o��4}Q(z�܄��F�gU�n��G�W���V��cJ�QF�8;��Yʋ���$���o��;�k%�*Cq�,� N�˘FkX'�ʊ�� ]	�fg�̏؇kPd|���.�ٟ�5�V��yEͷY�4p�O}����@�Q��<�3�Fy���~!w5�������׸>�4�:�˓~�#�|��D���3y!�o���5����~��#�蓀r{��k�-3�.NA���(��Hs�xԡ
*w��#U��_�i�h��O�N�]���\-y.D����\J?��b���z�b+���!@7����A��-QL��G-�{���n����rhX15�e&�K�U%[P1E�Tf�R���[��*q���Q�$ �E��:��n4Ca#�wvb���-���e	�wS�I#�%N�����!Im��������ͭ����G��&Z��0��]�'C��h/�� Ս�'��s�5��U
 AHQZ�H䌬���m���˝U�!.��Z��u��s��y�1�`�(��e����CL���뉌$�G��\��G�t�����ڑ��m	�6�&).yά�-A	YT�F�8��$��d��I4���&�Q��3	^(Z�Ye[�����0�4���L�C\�H�)���,0S�w�g�r|��r�i����C���?9뉜�!*�p]�[��۝z���h$AY�')9\�`��0u��b ��U���
A��<zۗf���n�n���ة�-�6Q��Cܵ5�!e���C'=O�Bo�6�����Oq��h��+%�f��x������H�;}����h����|>Zw�"l!C�7G%$��޶ì����&>�e��s#��\��6�G�)`J2PO�*iİ���#�������i�ճ���!��QZb(_΍��9���Ĉ&�3�0:��9�v
���uNXdP�m/�^��>����)�&Ǥᄆc���}�S�/�L�"O)O����`oC�v6;v�.��CH��.���|坻R���i�IV�E��1ʗ�6�������}��0i�my�!

E2a<n����s6J�V:����k�yِlnx#;��?<]��m�Y�2Uؒ\���Eތ�;�w#h��3,�j.�J!1���j�ˑ���e���o�;Gt�>RGq�"�O[3��2�6�_z�pG�9I5�S�G�6V	?l�&A��Xi�tItm�H�F3T��3r6{J#��#C��^e�?��I�f�Z�O~,�B��T�"����{���uM�f5a���Q=kDx������ �C��wg�/����;y���J	4�K����7�i_q�U�/��2ۓL��*@�e����T��ߺ7[_�W���)?��J�g|����QQ���QN~�]��l���e.GrJYc :h��쀢�K;߯�n��uBsa���E�'���8���!y�(��?���7����H#���Q���̋ռ`�2�}�e�@���8���}�	�A�t�⏣Q\֏�UNҽ�*��9��UqI��At�$�*p�o!�CeZ��R��}��GZ�\���!�����da��B�0#� �;G�G�Y��t[�����݃n��]��$��w���������[5���s���O��{�A�����]��t�c�,���}��Fi���Vó4m6��o����>�>t�	��P�D��P�8,e�Ǌe��l���&	#~<���~��.RE�Ʒ�M�@8�A^�g�͞��َ�_�J[3������J�:�ڝ᯾��p�3����%o�"e :x«�ҹ	~�	��$�t�N��_5�VJ/��@l���yHk�rd���@��K���g�C��}5��j�7z7Dr��G�!�h��q ��hd��JC��!+���+�}׆?���𚜍Fr&�b�J<�/�(,��gk��SA{�&�"��o���m/\C���8��KWF�!x��?aϰX����K��{k�t��C�1�Ô'�X�8Ø3���F4h�Ҁ��%��,_����G��YqK�^�Ec�qψ�"MG#B��1��F�.��qJ�0��b0,�{b�b�؁�ޜ���@
�u��������b�oe�$J�c�aJ��h�}͸v�V�[�ђ>���l.�V���s�p} �]L���M�&�����K�"k�-���"�m��%��M���.�����Y�>2%DEpZ(=�&��	O
��[��Q�� o����*�,�A���S��|��r�x��^�3��E��Rl��u*��j�G�'���6�w�����b?�on���nT.��*�Se.Ù��Ts�pD��J&�݊Y) ��'ur@v8��T
��X�Y6Y.����!DU1H :�V~ *o�)�����C�O�T�l:Eel=��>�����η���_�)����'��?�+]ZFMuf �KKb��y��71[�U��,c��j�����[��-Y���6� ��ر��c�w>k��Үo��Z$2g�(GGM��s+
,��%�2����P�\x:���ߢ(��#X�宝[�u-b|�6W�5��l��0�Z94����&u�M4�yj������q���$����-�5���;��w��"�>���e��
%����glQ���ܼ+��� �ә�K$I�f��K���Ġ�Y�$�ٿ9:��t��h<s�z��>���Y�.X"Q���F4�q���+�m&���V<����{	�''�=����@b&�L`c�	*t<����3G��	]\��j>+6�h`*s\* ~�;�E���-�0涗~_g{54���K�0G�U�bx!����s:(}D��J���]�X+��e��h!�"ǂ��?����.�C~\dO�W�s6�A�X?y� �<7j�a�:N�/�6��͹z)�����~E^�j�VhDqH����_��m���&̶��(���T���L�.. d�ʛ��Lw+2_�B�kA#�Si�s�f���E��_6�b	{}^%"�[�ȃ�X!1�������z�S ے.����)y���>��T��S����j���vM��+^)�f��z�D^�B�YV~j�/���r��W�fG�L��c�z'j�| D�.w\5�-%Ν���@��G�1��6��;�Gn�S��y<�08#�y��"���C.�n�5QY��RS�" iwkL�c0�e��J#��7@�
�ɏVn�w�a#�����(�#
d0�y���g�NR:8����Z�@��=� ��y�����T���V�x�Ǔn�21�
̿���o�1^l���9�����`sυ������y�M��yڰY�L�L���IL��Tl�I44`��*�6k�oTb�*):.���N��=�	*#;��C{M�q$	�ؘ�^e�#\#L�OY�*���u�Q[?p��w�o[<� R�e����3
ZL^`U�`a�H��{I<�C���=�G.�N;.������?��yP��j�<�r��e�}�;�[�KP1'X�I��M�� z���r$ދ759L�w_�	ĝ����*w�,���ȵ���t[C�C�C�1S�pg�D��b��m�r���w�&Ktd�{�w���Q��4�U7YJ��P�tv�գt��6Ax8�0�8��;��$AN	S�'1��&�1�$rQJdk웕7�#>u7������	�̙5_
O#��\�1��V�Z�n
ѹr.��q2�f^�RM+�"8y\�3,���'�,�k�Z㏹5�W%y�~���31��3�X�0�Jӳ.I��Q����fۊ�._I�T��B˄�C��-'���>|��7�L�*���R<g��B���%�0,��}�+O�j1$qQ�5��!y�2�uQx陭˙�S��^��zx�1!H�;����`10��T�ܗ��=�M�� vt�#�6��K���}�C�C�?� ��fu��V��$7[��T�4B�؆�`��F�!��e����$hN1�<���(3��G(�Df@��I'��b\q�!zr#I���CW���w%�Zݴ^jV�S�Ҕ �=�[�*	�����7��}~B�����՜��T́\�[�骞��w�f�-o7�4b�}<��	��W�3)�$�l�<��넷�*a��r��3XY�ճ؟]OdAm���\�'rˈ� ��;���E�Zo�LX݀Βlt���=n�Zu�%��l����4�q��ATH�9����kU��[J0�B����+'�(�:��έ6��ܳd)I����yN�|p�Yף ��&�]¿NX`|W��:��#�W��S�y��35J��ׄ�N�N�	���9^8�Q-�.`��l�mI���c��H>͔
S�.l���u�^��났|��{�yb��|�S��`��D8[=I�|(]j)qb��0B�)	�=R�]�1�;��<���?K>P�rt��
���l���0Y\����}�����[=Ek$����I�K�V�����Ԋ�8�J&0�8�?��o��<�I9dtm���t��$�8}-�8�$��'rC�4���gy�eb7=)��bB��b�lJ��a����V��w�go�;(��@���O��f��ӵ�Yt�4��n���?��9�5�L����O��P��R0(KB�h�):^�������1$����]7ٯP	��4A�S:-;4�1�ӣ,&�SVsD�>�D�YBG�p��N��ꑣv�v��ԕ���=��KlEc\|�b8{�қ�	���������V��9-x���������S,������d��a���8�v�<��Ð1m �F���{/�97���ADΐ�tX���ta��F%8�d�H;ȇ��EE��I����:'P,$�p�ߙS'w�̙�d
����D8� ��oc��v#���xn+�4���8�����y����?��C�x�<���1��5R�s�BZ��o�� ��E�B1�c|��mǌ{-p��Pע]�]P�y���l����u>C%c��Ꭷ��nx�?^i`;�sR� �f�����Q��=�R�ȇQ�|��X����~�Y=�Qw���(�)	-�h�"2���*�2�W�3-����dƙ@=�oJ����������?VmUC<ngCSI(�)5?���Tp
�<G�1��/�L���wL�p`�G�XB-�� ���U�u�<�\4 M�\iiʗ�����&0	E¨n{=�S�!�Ƃŉt��0�+��	v�@��Ջ�7�S���YO�SG��𥯝}"�CAʧ!hd���Г��\^��BRP���;��mv ��\"��.1	��R���&ŝet띑zl��1N��*�N �Znr�:Gb��G�R�3���OȆ��Ŝ�<��\�#���x���@Vu��|No�_��?��6Ipu綆�=��G��R�?���M�˅�Oa���vp�/���q���,�@oM��K_�!?:��3�M�@(�CŃ֢1G-?Ci\2lS�P�"�G�SĈ���IAa,���6D�I_C�!b��ai`�#��\v�{Lr��ĖBAM�q�*lg�δy�3�[=(�R�N&��}���i^��� ��uղ)��I�/��fV�c����A�<;$%��*� ���+T"�xQ�'ڹ��y��Z}��o�풗D��C���/i��*���{K�٣�h��b�'��@�н�a�P���S)������o,�?(�
��풶T��Z�x�.@@��W!�e�ܽ&�\�R�(�uc	�q*E�1�`J�-P�nT�
��A����a^�@�z�#<��څ���3��<#��cRS�~�z��Pa�;��0�b�\�B-q����[�"��\���k}ϣ�IٰE+�<E&&j�:��}�7?D�� V����U�w-�E�!�^�-��8_��)��E���=�j^���FA�τB���֙�|���RUBOō��I����b�aB�q�>�iũ���)����g�u0��K\]]�}F5�[ �S�{�z�Ϡ
CN���|�2�����M3�<<����H��1��z`�{�`;���HMb�\a�]rj�Y�Y����ӄ?>/O�i�Э�+��������\��tM�a]{0Z�N�t_ �/"B}���s�TȟBt.ANΰ0�y��ku4�ͨY��T~����}�S��^!̧��7۩,����
4K{cc�5��9���������D���Bc�M��jf HVog�������@V���k���j{�����\�}�+}v��N�.���.��2{��b�*�:�UXDLS=Ѵ�K�(�	��|�άb�hU'��"���6G���[�Xh��� e��]@�AQ�}7����&q���+�)M��bW��ݦ�t��'x���5����054,*J�ޫ�X����-��+��Ct�{�2
�8y�J�U@�MI
�(��y��ag
�4D�:V������r�C����)�''�\�Ҍ���eqi�Ά��JRw��[%䉙�ՐMv��d��3��N�kc�y�Q�� �nƒgR-�/�TJ�і�W��\���=I!���}+�
sh0&�Xe=��2;J�h�"�d.ˮVi�L��HwcBq]�]Nl?�������z��$fD�I؆�5�&�DF��	cn{�"��<���9��4�)i"��#
��od�����7$��T�<��-�7�?q�ܤp�3y�3�I��#�wV�"n�}�����}���̑2�0�l��m*W����B��Q=h������YW�KhU�ğ'��.	!6�L�Yg��4D��h�
���i��6�i֡�p�����p�ة֒;�>���nɀ
��ߣ>~z[�<%��i8�!#�N4�*�n.Y�(�Gv�Fl�Ϗ��"=�M��M��oc�c��Mu2��";G�/v
T��+qn=#)���q�I��7*9࣢���/�����rZN��]?�l� �R��f�8�֊6�a#(PN�p»к��k�����XN�GQ���`��!�֩x���a����M�Q_���zwG^��8�Y����5�fOBv4��/!�Qݟ�-g~�?���M9 ,"`"=�)e�S�뱙��d��{͸��Iem�q���Fz��ڟ��N}�?����
^�R��1�/ѭ6C2��f1�):W�1-�(�+��|����G��sU�X��XVA1D%�x�w�eP�����],#��5����P�pm(�Տ���?U-tꗪL<:�st_����n��j��عR�Y�����]��c���!����Y��b���e��4&�˥��E�T�I���ʀ; ��x,�띹9��@��Zs�u/�H�G��Z�v�.�Ķ���8/"��S�r\���笭�w���}�N�}K�?~�������^����u�"왷��d���{C�v�k�C���IS��y�4�������|��i^�i�m`�aH����l�p��DC������$ć�k��g�EZ|�h$b��ƨ!A�l�U��ּ2�"���<���S9&��O��X��g�a���%�D�e��L�
�f����-�:+�-��_��J/ $�W>�j S����F��eI뾜�J�-/�2��1��f�[�L�-�f�{A������ƴ
,�}�Y�2�QZƎ��&�g�5(�\(ь�} �p?+�k��\@� |@B)���A	 8�@1N>Ҕj����گ�X��me���(�E�r�Ҍ��{��Rc��7�~�	�JI�����7�k��=��g�&��f QDŇ7{��@z0Jt�\�Y�6�9�Z����|�o�w"��IY���[���|��^��E]�_���"��T%ZZ����O��|X26g��w�b���#�Ϟ�]�s�޸��:zӓ©q�y��_[rHW��û杆Nt@���=h�ηN/�}A��kk>P�l�q��\.<-�%��)k��N�*xOϝ	
sz�1��=<lR��,mޅ��\��9�g�|��v�0�|S�գi��eO��Ù:~?�1�j1�6{�g��ځ��8E��'U�$J�4��$g��˱�ܸ�A�d�/���xʄ�N�{��>�{��"фx灎�8t��vS���?�q�A�AbY�i��")C�q�/�V���=�Y�� �R���q���j�ެ�j[Wm� ��<��- ,Co��4��v�}TCP�-ʞ�Ɖ�V�q�[=��&���I��J�H�����;?y"C�йU�-�<���	������ɡO�������i��}����B.�o�b���
Ń�R�r�4B?6�M}`Ir�0J�9|���y)M�q�.yZ��能J{�\��)y}�/�T��������,)�F�Y�X@�f5��y��tz>k;-5��a�6����.�gc�	��˴���}κ~�.˺��*��=�j�ᶡ��������Z�3��]x]�u���v�wVGjĽ���R��h�5�Z�x\�%����A6Z��m�����
���V��3]w�"K�&�c�v�T�wE�Ek��6۝Jt�H)0���6H�B���.b�-���Xp�^ˊ�$Ō�Zg ���n����(�/w���hѴs�Co�	|��"��6{T��7�)�e-n����1oZ���E��M��|Z+۞�J�ܨYQQ-3rO
s5+��i*M#�f��U���5�M�Q�S�EJ]�C�:��c�d��i��-���Z%�(�:t�ok-��/G9�iw�P?T�9 �!zX��C�Q��K�G�Sr���3
������|���y�v;��=�u��7�Q����Nc�@UWP���`�6-o�68>������q�y(���q�����902�f�"`�:�i�BOdz+���JvC-X��m)�x�ņ%����ɯv(O��n�-|���n������+d��#�
�n�b���4M�r��Ƅ8�S{�u
؀�)!§��1�vLvY�uOS���}�v(��bM$G�����Z��h��:�kڅ�We�R*�2�	��q�>�e������3�ia�})w۸�z�Ā�_���N�D�(W�/�j��||Q���H��@3�Su.(2�0���e�I�n�nD���K�^�z� ���Z��8p����|��64�}���ٴy�B��� ��'㈬<���w�4�����7��co�-�ŷ�y� 1��$��$ǯd�K�����)�+ �u�"��)R��ڞu��;��oY�v!�Fגv�k�7�Z�	$�d���FYwL�A�ጛߣ�g�D�|=�ԔJ}C�T��?�"�'_� ��	�=*\��H	&-��"z������?����#�e�6��=Օw�T�4�u�����Q���t��Ӈ�\ҹ�_hg-6B'M�2��D+��\s��
�4�!6�/�(�nN �����6-4�"1�o�:'b��.=���p�,�.ô���ѿ����D��1�3P��G�Ro$ܱO풛��d~�'+=��~�	��Cd���;� ��� ��ũ��cN>����{�]����Ų5M��7�X���EU�NιҦԇ#��Pt�w�7�������Л��'�V��S����_�P`�����(���!dr���Ёܚ<#�.���E��P�h\����2ٳ
�	8�F���n����}O;�.\�6T:3��0���}�%k�~�� �3DA0��j��q���R��2{;H�)��v'��c6Y���� ��G����:�W�«�t,&�)�
�a(j�>b~�F����@x��1��`�y��O�S���~�cd٦�ףּ��tCh���fտ�<���@J6��C��ATu�M��(J�t�#��LS_`���joS�L�L$���}�Ԁ�*_j���0�	q�)K��qu��B+���웻�f{�֏�>H��$M����F�?�;>��4�����`�-3�3�X��p=1G��y�� �nw���/�$\����]xd\|������_Rrm���6P@�h��7�6�/27�?G-p?�S�F�3c|	�_�b��Z��Z������+���x�3�Ryfj�:�� �HD/{�Ж����/3�	އpm�aW��m�"S��1��pe��lxyǚSb����_�g%POS�PN�W�R�ZCc�
Z/�+���qB����jD��0����$;�Qq��pYs(�����p'��eN|�YM�=�=��N������Ԅ�Z2a�~�"����N�+E�����?G����;1���n�k���0ӟ0L�jl�[��$�����P� ?�S>�:�*f�k#e^���l�W=rZ�z���=��_�J���[�ىKN��Z/R׶�mٌ�{G)*���i�˗N�/��\ƇuJZL_������ZX��=�y�������H����Āw�:�!m���},�V�Æ:֓]��֢���	d���/��$�n@*���޹Yc���E�6���.`���u�ɩh= e�]�6�O�j���g*o�5�!J��?\��bS����*�u��!E�s��"v�AE�_�������wf�ג��
��8_)���Sb)�0rRq����5t[RL�fTgJ�ڏ����Rvj=�AHv�8���tX�T&�+TG�
�-.�˵��$� ޝĆC���yt��w��)u�щ�WWs(jƠ����:p�K�Q��8! ��]��m��/ �ӧ�L���������N/�n0~\��l=�s��=�ԁ��@�$i��Je��X�!�}D����	z�Ѫ��[q̜��[T���K�$�*GVy��������׎mnL�1ܑ�8(�apYu^"��fI���*y@�M���Z�-���ݾ�Ō#?��J�񩂠v�ڧ<�!W��STPo~)g/��!�c,�����6���{��u-�5%���a1f�����Q��Nr��Ê�#�X�̽=��䯏&�znb�9�>��?nGjȁ�sm�[�v	��|	�;�R�H�Gܑ)&�?���$���쌳2'b��ℌ��5��f�ף��{@��=��z�2dG�魛7��0H��L�p=u8�>����0�q5&O��;X�
-�daM���}՞zUo�A�5���0�>�#|�:'�I��T!\�1�"À`J;�̖ov�/�)���X����v�kϰ{�yV�*L��*1~.\G꿝�������\��m�;��m𲱍\�V���������}Jwޤ�s�l��=ed��W>��w �M�e�&� ��`i�6�����dG3;��`�4	����_[���wg��q���?R���Wcc�F����p4����k~��
��>�OX�b�#ו�4�c߯�C�����.�Uʍ�ƻ���%����偝��A%�d�j�r|���ȱ�^�����ie�'�����;%�}���{p~m$ ��
�ug+��S���x� �Ԍ3E�+�=�:��J��1���!��D�'�M?Mz[ZeS�՗U)/ T��o�85V_fO���h� ������J�ϥ2p�-�i�@"�`\��2��l���x�f���
�qb�A� ��}���1@o�u���j�W�[C:�봢��]v�M�8�2.َx4E��``
w��賯���1��W��Hkf����"�8Vm'��ا�HVVI���6���g��롬D�_嵢A�Gﺴſ<~�r��^e!�~ȑ��H��g��*�����a*Z4	G� �� �(����?Ὂ�������~!��=�6~kQ5}K���
V�t8$��u\�l8��.`([J���a�5����>�{���^Ȉ��`y�8d��P��^uP5���s6
�f���w�f����W�"^�c�}�;��N�ɺ�L��f���7%��1��H%�W�'��� `�=4�����H���|
p�v��ld;���K�ƥD����E��M� �G����UD��s��!�6f�ϭ�7᫘������Z�Y�8�g%n�^؉��}3�Zh5�Zظ7�տɖ/�潪��݁��{�Q4�>6�n���\;o#�L
�{5��n�j������	����<�顆gy�����-�Q�Rl,��$��9�"j��I�D�ȳ+���<������J��II`���Xr�C�%[.|i���pvDcn�=7�*�2e��V����J�G�l$}����f�9DN�Qв�����c.Lf�4t���<.Y�!�ɱ�ٰ�;�|B��7�Ѩ�xB���9��oڱ������R��e2�V��FmW �Z	p���ЙIO+���������ߦed�rCN 5���%�%��S�V,u�P|kK��&O�iO��+7������D�g�����4-�L�>VA5O���+�z�9F7����`�E�3U��m�[��R@��&O:��v0��/��G+��#bj������B{��NC���ʯ�b��N���j`u����q؆����_n�D������5�	���k��(�Ys�XKY=��u��*SK�W�Rq�����^�G=�D��)�~�rɺ�aME�:���95ᔜ��&8E 1T�z |���CB�o#�y�m%��3��� ,��ԫւg^��E�����Vn�XU�|�F���O�DԻ�J&� ��E9Q�"�2����w�Ȟ'�q��$�F�����=;����E���̠��B��,�>\���^��y'���:\\x�a��E��{�n�j��35��=J�_���:����ԾS��s���^�E��ΔcU^ی�Y�������_�����3߮�z�#`T�P�b�?xx���_aeQd�K�AvlA��x�:�1�(��E���"4�Mo��0o�hh$�������t>��s+�Wz���Ǔ=�HGaqИ�n���N�'�YqT,���k�.�ڧ���$�~f�~n���uo�(|y|�E�0�� �Px��q"ƶv�������&��'�(ɸ�zd8���4�%�[���B����@���Ft2�n0r4�>I?��H7�GN.L�A>Cv�=���Ĺ_���$ ̮�"j��ǹ+P;l?c\�͙���8c�����ahԢ���B��1���i�����	���m���H]Vp������s�DnxOܚX�Fb@��!1G�gb���e�|�;Snh/)�\yS��Ԟ��<��p���#�M�XH>+���i��4�� ���J�z�vvj�ײ�|^�g֘C"TA�Y��C@�[a�|�kG��n����ȿV}���fh��o�_̅l���wU~���;�+˖E�/G��W��6���LAr� �:)����+z�j ��5�n�V���hXE�;O��:q��*1�4�
!]�AQG�|�^�n"���8Y�A�%k�0B˷�Qժ:�m��V@@�O��Ԡ�]���Τ��m�Q�r[p��䏭�#6'� 1����-I���[۟��{U?*��a���*x��#��$rzCy|�����2���m@�M�}��
>	X�7(t�/2��Wa��,}�^ߺׁ���0E
ƒ0huڳ�:MW	�$G��*�ē�_��羍ۈt�[��x�7�79F��$�����t�]E.����� �V�u�oYm1~Uj�|�w<6= 4Ƭ�&�jUA�z3������R[�Ŧ���0F�!�f���63�z���C���WD][��Z���(6��v�"�y*�-��Jaj�'�ο.~�{��W��O��o�M�P�8=�<���s����m��rܘ�?P�2��wX��Hyki L�Z �ɒ��9�O�)�-j�T���,��Z$�ұ�����^_�\MZmUs�(6t�HX��H�sEŘ�TTQWz�-sk�w���l�L�\*��]7�}]z������|U�k�`#O�2��O����e��YѦZ�$0�Wtv�$� $�e|e��$L�!%r�R?&h#�+�@���<Yj\�;�"Ao�0�K.0NZ�]��YvP�!R)�qk �,�D/�G:�兺�@�>]k��&(�"��ּ��^��T�ͬ���~�.�P�IQ�B������f3���]�`��b~�Y�{@ ynA���R�{.���f�:o�5�{DW�{�'b|��<6z �<$���js9�[�I�}N~ࡿ{��M�3 ����ek���+���T����'�bˋG��]��	;���3��0>��v}��6g���N�K��t-Ϧt�6X�]68�ɶN��Q�p~��5{(��r��p/{ ���>��P�0[��?Bk�"�Nu���S��2�-��yS������q�������u�Y8��]]:��ta�ŜA�z�8'��*F��!���Y3L��~��m�E0���I��@��M�WZ�I@=8�w᜸��-C7��h��8E��x�G���7)]�~�����+�����OO�����yO�:sM���㺖:a7���e�������V���1�j�}��ģ�4�:pG�X�����֯x���dm����՝d�k�MA�5�W�o+�x�	�
�����H0�c�ǫ�I�wȇ�` �i�0�,�z�\�9hE� ��C�S��^4z9� ��o��.�N|>gS��3���[�D��zh�������9կ��>�&�c"�G:����g�a�����K��dd�"?zbf��+	WW*m����Kl��%sr^Ëk�l�L	��m�����N�d--uRHo�U��cd�UtYB�6��$.u�h�"�W���N�R5g$B�l�j	� �Iq���:���(�p8\�Ol�ԕJ x-'��H�h����!W���JN�E�Y��bMD2ⲩ��%qA���fWɵ�x��~R`�Ծ��`��\6��D��(#���\�X,C48�v�10��i���X������`ʀ�X�Mc]����B5	�E W곾m�-���j`�͒�j�g�:�_�\����;����	�V#n$z4 �Kӂ����o���F\b������ѣXdp>���ؓ�E�%&�d���h�,`��	8��U����Ϸ�� e�c�����|:VRXx��O$�u�s��%�Θh+�)~JA��Ș�'���d�����a��w�\��A�����q��Z,�o��.Ǚ��BSO��$x'�hp8����.I�Fk<s?z6�@iB��}Y)�K�ʜt����B"��Pq�#h����qx-8�XA�`}o8�(D���N����E9���_�p��iZ�5ɲ�1��8���<y2�3b.!��I:G�#8IyԺ�6:ﺬiǪ��h��m������+�������Tν��ש�(��3�+(�a�l��ۛ�g����G�_��Y��.��M"#!��p����0j�?v����)����m/��J:�w٣7��?J~c:�z��;�Mѻ���=��̮Rm�k���lֶ�v����-�!�z��i�a��6cZ_DX�*��ݧt��h��Jc���[a���]�1%���;W���rd���1�F����<�¸��Cn+y}��?�T��~kA
�#��@��O�؛9|^Q�0}�H>��?pL��jq�t@���/����w^��>�swRu�C&L3tΕ3-]�@���_D;U���HH��Ƭ회FV���rau�e4}���:�Lѧt`H�s�(����)ǐ�Ԅ��=�=��O����O�����嚄�"�"T5e�0��#�}=xI�"~Ϥ$��Xm6P�r�i��g��r���mS��c;�Qq������������ч
z�Y��ǚ�z�|�H�ᄀMkF��=k�N�x1�0B�
��x`�����C-O�XOBm� �u@�D��u��9��Y:���
{��"]aYr��i+�P���:���^�4Ky�/�n�/�C����W�������c��\3���_��w��.K��I߻t������#���Jh��V���!�0	��ช]QI�6�tvp��sЅ��v��������os�����.���o
o%��=f�F�yO�6��|�b�>#�U�^J��3�4�E÷'zV�LU+����a�,R�裌���@�s����������:u����|����}h+�)����M���^r>��Rj�8�?�ʜnc"1�/�=�^�Y��S�j�U,���k��܎$&+�L�5��vl�{��0�̯�j��� �W/U(��VJ�?�76�t���m�BJ���sn0������S9��ۘ�U�]*�5�^}�e� Q�X��	�J�6�j�������-��
>)k;D&W����ۄ���L�}
��M��_	b㉳b���]�ܚ}��b�GqS�k(��_\��5y"��0�d߻������Ear���K1�$F;,y{o}�u����K�k�{:���^b&����8�o�r��qq���;Zz��@t�4U�^:�?�Q��/��TՋ9�Z��$�@�*ޠ;<qA��QECB�f��N�8��� ���};�W<�h�f��Uv�C�m�F7�Y��/�C�-�"ߡ���u��.�8K�c�i���6/�z��Y���z��q445^�5!_��=�,�wR�{#�������D�)����r�}[��y�
� g���+I<�D�9�jo�!�4�D�X�3�����{��W��M�	�x�ф����+��&S�Ҿzv�ך���U̽1_�)��P!���sd��L������
�y�=m�k@�;���ᝬ�?l��C-�DC�D�3�Y��N��v6g~�O�vU���]�|O�|����ocJK0��;NH���������N�P���.���5��NV��+P�0�%h~yj��@*���BI�WW_
��Bț�׳�B2�1p�e;5�����6kу�'�!F���bI���Ω���yj�[z�%��*cN
19f�7&g�����%Eg�l�ކ�W��w��Tr�&B.R�R0�1֔�\�jZޞ��u�]�O�"�;ԡ��|���_W�"��� C���j�l�kʑB��p�i1=c$Ib���Uih��"�S��W̳�8o�lfj&�<	I�ˣ%�94(�k������+�V	�5�Z��Q#�̍o�Me1��w��ˠ��jvIC�W���$F�aZUV�0P��nl���Hp#���_�A����Xj�}����f���5Q��h9�ii��G=¬���f�R��lP�=v6����V4�7�>���.���/��sa���r��~xh$$��~��h hCQ�<ܽFp�y���!~pٜ��Fp�8���y�6wsY1q͊�o#��U}�`�9E9f_���F��y]aT6y���L59�g�fep�+A�~|��2�-�j����آcd��W�����g�>Z7bG���?2�hr�N��_|�9.s��c{�ho�__�Y��}���˙�Y"N�d��G�ȱ
��]>�'Y��0@9�o��R�kYz~��P�A|Td(�	X�oz������A0��.���̓��QlU��H�+g\�j����%�Х��r"]%1����Rq�����S&_/� f�,��]���X�1��ϓ���qD~���a���˻!&�|�1��)�n��e��R������^�u���<��5� b��d�Hk�+�3�h�f8/�øB�N�9X�੺8��a�Ɉ���;�����q|��Q֮ۃ��j���?ʶ�����-����{�X�
x�y�أ���5y���+��Y��P�*/�.f��a���:+�VB��Ĉ�[WV��/f:D�c�.�M�x6�FXe��Zˀ��,۪�K��r�2��Q�5dAx����ޏoo��^��n�I|�MfC�z�v��"�����<z|9��N���ڟNr;�9���I�*e���f�-M�N,�T��&÷p����K
TD��������	���et�A���S�R�+�, �+e�cCS�]���?��P�Г[6β?����|<�C���E`h�\�f�7�T��/����/'��g�D�Ѕ�*U3����,�r�ݪH1'|�<��IM�k,Y2h������'h*�Dm�f!�aY0 ��ᮒ�������.�����4����,J��/C&z�j��mڍ~��m�W֞߁���v�zF�[������z���K9��	1��������S��"��.vz.^�RH,o)v������7]d�5�nTUQ��٬�]R7Ä@��/m�yt�9�7�w��7v�����x��v�/�W�tV[����'7>=vO���UE��5�,A���������������tpw�	��p�o��?�ˬi�:U��>Uݦ,��%$� �ս��.�6�߾��Y�vG����1�����	K��@��w��#�gR
��Z�Ze���e\�=��@���rڋ�w��]��U�#�㗯���%0��f�$�����������X`�Z���<��Ri?�
��k��%�)��޼$rP��o]U�l-Y�e����jޥ�)&�c�n����������Wfqi��P����������Ǔ�k�<젭������B"Bb8��+o�*���2�K��o�c��p�"�UB�'��ͳ�W5�K�F�8̲p[`��2j�Ȟ�M����D�ێ@�y�v�Ӗ�T�re�{Ϥ��,#�xi�K�������#�k~A�p	�Le��}ŗ�_ZW:��sO|�(�s�c��Z����48�~��뻉�K o��>I�˴�\Ai��5��1y$P� ^ĸ�}v_�Y�Q<�BoK�A�:N�����ƶ�Ǌ�"���u�����$�W�W��:N
Ў�E"˿�_u[�<�4#d��G��	>�����U+���:�'SK
Z_��9���2~?K�j*/��u�u�ᔝ­�V$Ǐ�5���ᵵI�z�|Y^X��T�w�5�h{i;�j��Z_���X`�L{��\5��M#WҐL�O]rz�/E��g����k*5r�]���l��7i_����'���T��w�H�u�>�pu.���!�X���yN�u$�X������38�}���g�W�s$��0\M{P�d-o�n?&�~(����䞆�S��[G�%�òSV���g�3;
$�`��o��|)��@ʨ���7i�,QJF�giYr�:OH`ǻ8�2�ݟo�l����@S9��͓�#RH���+󝽻�����=O�~�f�"��_ZZ��.����b��o�|�	�y5\__���+���7#>ZNr�H�U��5���}��׬ll�9���U0ddAdτL��K�{��,��`c
��E`h?���NЉ��Q��_>D�
�W���78����U�ЭF�J�FwA��OՓ}�`��	�EM�N��H��&CD}K[�f�D�ySMMM��@B�q{�kzİ�gԬ����?,�*A�������vt�v?���+=]����jF��l������Ieh�BV2��6`������Owg�@�N��Z��������v�����p��r��Dv<�2��p�������)�ھ��S��m��႘ѐ�"A��210/��"ً& ?��1��zZ�Q|�����	S�����l~�sg�ٶj�K;o�j�ׯ_(5E�PC��a۶]iX�k)����`���i���qi�f���,v�����pB�s�EFO��顸L-��v%���Ƅ�������vQ^�s5�Hu1����t�;\�*��۱�u�@������;����XԨT��z�'{����dM/L��*mq8F����/F��F���C����٩GQ��j��i�%��n��`gar��4O�|�p��a�?�CY9���a	_B^��?���<lщs��upa��E�w�~x
��2�\9\:�
�=�=���e�nĄ��#TӶ>"F5�DLx�ؒ^�F���j�B �7�Ǳ_�������Q��[��Z��7�zg�zn]��G����S�i!'�b}���ژN�/-E�l�+S�KYN��f�ށ��L? |��p]ؽ�5��Z̠�e�ҁN��L?β�q��=�����A���=�w���p��z���*���C@K�ww�T�P��V��y��fٚ�B;�9��r�h�����?�z{)��,�8.�q�\d�R"��8�� ՘���ݢ��Rz��t�����X�v\��
h�V�IP��	� �T��g�u,��p�NM݋�u�I�ĳ�׌S]96��c:zٚmh�*�
��I���m�I��N�@NE�����Ŭ���p���>�B���@������j�O�����P��ݝ��ۛ!N�FJz*�'	��=��܊�}�=��=;�X�������Z��
lG�i��h�"�m`�K;�c+Oɒ��T.$�^���h�b[��z���d���;&����d����G�.l��"h�=�`��y��8h}�� |�V4P)JG��pQ���ZD���`��=Hɔ�����A��2
r�?@�i�."s�'b�6���哟S�o~�u���ʻwEH�4��|y�H�l���#?�3m^]]�DF��1��\��d%�����;�L�|��C��{V���8S(�4����BП�����|���
�:�ల���J�����剽0֍*Xwe����V
���,[�UW;�e}lX�,�x����(~��sh?�O�?ȧ8B����^$V��ga���-��ɉU�Dt�c�CKU�����eTW������^��p�鿩�#��2bUbkn�z�ps���5ဥ͉}��S��!��u�~�� (��A��ڪ�w|�(�ϩ�&R0$����'��A�r�{Yjp �p+(KD�^Y;ձy�.���q�6����'�j�zT�Y�ɜ�M� p������[y��Ĥx�/�� r�F��JeKC�J�m)���=n��6i`�'b��4]� J_���su,о{�����Fy���Yb�R���o(a�-��n��V���w`�����{\Es;Ι<o�ܝ�Ue�z|� �=sqe�%��m;����x��/��o��^�3�e}��Z���xSEu�ZQ���)̎�F_�p��-i֯8��hռ.k ]��6Jw��	Ҽ��� w
U���:;h��-:Lk�c�."�:���M�e��z�9C����v�[ׂ����l��UQt�ID���U�(e������VGc��c��:	�����u-&��)���ķ��U"�����?�ϲA���ө�;�i`��#}�V �ic��a��RG�li!@Lq�<�a��)��˽Ǉ��`H�L��(�O
JY��-���R��Y�GTs� YFﲭz�՗�EqFbZ'��� ��y���FE� �@��A���L�����E�?�$��F����-kQڨdK�ik߁C�����N̳��k_(6����P|ּ�������X�l(<���iW��K�D��r�BRIו]WV����ȶ���Z�4bU��Ѩٕ���T�9Z%3���N=l�P� �_YOZ�t��>�%+C�Q� ���ɿq�7����� ���vC��8b��<�#}�9b>�/��B�o���bM�<P��@R�E�z�{FN1��z�0Ҁ���*�[
'	"3{�v3���n����co�
�+,A�`+����>ͱC��RH.i1|��V�d,3�3�\o�4EiU2 �p	��g�n�"J$��9R{k8pQ,h���fP�
t"����~	 %��y2�f���G\�r~Ј'�{�RNF����NNC��[���C�����AW������g
�s�V-���0����(<zAh�e����,4"g�돡�&�A�L8J���"ĥT��SNQ%��$9���1B^tdVy�O��t(��ϛ���Jj���ԭ��~C�R��L:�A
��gI�`ޏ:�Ҡ���u����*���O萹�B��8�0,:9r������p�U�*Ñ��P���΢���\��
���n��=U�@�B�Fk���Jy'��%����g�֟�dj�u�?㻃�p�����+��lM&z����Q<�Wrg˗Wؖ�c������=���qA},���fKqdEO��?�o��ԐR>$?6�y�4q������`�	���x���n�ʾU7�t`�Ă�X�| �B�åE{����������`Y��xVV�Q����}�Z�4S��D.?�ztg�j{`_�J�죝�O�K.�����o:�D	2^:�S��(�'ws���A�O':P_<���[�ŪY���{��q>	�<��L[�m�e<_��Ta.'2x���]7*�#�`�9 �z*e��!�!��WY�x�u�x���?	������.�ZА>^�r7����~��Y�c�a�$H�5Ԯ�f�$��vԜ.��ݺ	�0B��kZ��������pX���sG����g�$7�H�jPN��@�d8�q@ۏ$~�����^�߬�k��擡�H:�Љr�m:��ܚ]:W�b�?�r�D�T͔�HFބi�}>G����3�`f�p�΀��|lϑ�LEʶ7�:�#���gF��{���WW?c%�!�`i��fk �pD)�g�7�vN	A�Ә���ʼ}��>��ސ��I���8�AiW�lF8f�:�?b3�)�����+\�o�Y�/J���K�����ja������3�_'��}c�
1,}��ٛ*�vvy��^J0Z �~��/vC�yT�ck��:�;��bgU�[����	G���!�����%�:�p1���YK�d{�A2oG
��r�d&H>HyD�(p�re�h�d�B,s�I
n���BL! �Vg�V�p"�}cu���;�[�;`�#+|�L3L�(��oǰ۫��T ?K�um�� ��Hu���<q�f3z��O K�z����6��D�U�ۘ�����G��v'u�y����2Mo�i��*`J�a%�a93�����g+��Է\k�t�Q-��&�C�@�0L�hxgV,F���%}|�g��ۮ����ތ���FU��J�`H������|���߼��nܶ~ytd�s�7s^��e���"?����I�IT�+���;�[�Da���M�V�D{���ٕ��Ü�]/1~|'�4�o#.�={��;M�õl~�����6^���A�A�=����A�Й�ɽTuS!��O�
G��^U9ri� �6�F�K��E��]9a&��~�hz����9�r��l��¿"^�����l����N*Dv}��� ��>�L�z���o�� ڪ�Q�CFcJtu�)���o�\alDtY��݂Q�<��N_���]���@+�2x�`�a9Z!�ehT��4�\G��}����>�AFY3h�{�?k!*|�[�v�n��-1R�u�A��$��#�`����m��|�[h��I�ϪpX�VT��#L=F=p�ec�r�M`�����(8=7��2^�8m�`��|m�!\g��9K����l�|`�F�n羟���W	�|J�K��ws-�`Q�X�E��s�!��c;��9��j���(t���8S������_��Y��]�^B���FQ������Mգ��4˘��,�?�� FCL���~�~L�ň�ѡ��a�� ������vZU�ͮ���Ꙉm��m!�"+g# ���K�;��2<�C��ryQ=�D�%6�Y^����4Q� b!�)��K��L�T6ւ� ��4�)��n���lv�i?�x����0/sd05t����X&����������=E��TF7u���7%܎N�J�z��IZJ{Xߴ ��z�l�=3X(���:{�9Mh�l#�1�9n��^�1y�Ȑ�-��LA*p���fO\�{�0�]*��~�{�EA�q)�b�vU��~��{��p^��r���1�����ŰF*��T毓��o�z���q��9�<��}�BN�80�Q(<Ì�`��5N����y9ٳ_+�|_�x��^��x8�C�fU�[������%@)�C^4o��fmcUOl�ݟy�H�#CS���$lî}�s��_�$]2�A����ٲ���]�Z�bQ�U�d��6B���Q�9"V>/}��G��$��QRp=�
�hR�#L
K���m'ʺ/��	_Ic�YH1^0��	��7ġ^� �g���y���S �h��'�$s�]/���G۾���HJq��s/t}l�5����[;}6��s_��K��{8�������@"j:��{r�LC�<�j��3�th�U���<!���2˯�o�vx�_B����澾:Q�\7g�3�� �R���^7U<�M�	O�N����
�s�V�aB.u�S�Eg�ٺ���%�0���2���wbuppQ��J?,�!��3�N|�M��1���(T����8�����<bzj��H.T't��*�@�|��O =a�0ꃃX��zw�&�2�Lez3��U�e���]����a#�ɳ�)��`<�z�lT,��Q�	M���ĲPƻV��EG��	�i�6�As�rM�ؖ	��2�Ĵ���܇ύ���*S�h+� ��FS�"�C�:�8?&�;��'T�;����i��V�u�̩�bM��������,�^N^�8�ǜ��hl�������:\'�b����h�ҡ��i�
���\�h�ޗgi'<m?�G���*�L��8�d��1�����
���Q�r��K>�/��s����x��~�@3��A4̽J�)��p\}.*�W=������Qh(��).L��ͦy�8y�X�E�fjM=2-����g+���k��D
Z�.��ʌ2���ܰ'3l��A��	l� �8mq_����\-L4����{�����\���g��`[�~�W堳w6A~����`7�ؼszړw/��[�0i7QC���谙S9�0�ҝc�1Ԩ�:S��?�;9��F�����=#b�ו"VG'z�-V�V$r����7�r<�JT��z��}	%_hy�-�O�����̓@�`INk��K�\��.9�b�:�x
�r�]�5�ӼW���`6�i�p?&����r��EAR�e����p����
�0�7��R�ۋ�4Z�/�C��lܿ��c��%5u{��knq��LB��j�f�g����o��꾰~#�^��.1Z���ѯ۩�yv�r4�2����|���R~u�=����
��py����lY~�1S�0sW�%�@p���*a�dT�s������L�`tX�77eFEC�Xuڽ6��?`:0Hf�׺���@}����[=*�X���a�&E�ygi�V��i�Ix��t�_�-�|��@��]5��\��?UaB�h�6��N]��� ڛ%4��YJ�i϶�ð�mkT>Yy<���?��S0"\�o�E+`��j*�p���PG��y�W���k��n�A2\�����
&i�Ry�D�ԕ1��`�!��)&9��x!'R@���A"5I� �������[����z��#|q�>zO�����˧�Pj���I��C�g�;8�P����$��b�- Y�%峲��E\-9��|�і
mA�n�@�v
EjㇻZ��M У�����y)%$�V,*.�1��҆F��E��ms��7"Y[O��!EԜ멑r�߯/�:�v���F�|�����r/�������z�T���5R9D�<4v������c܂hp_X8'l�>  �8Ld�&���b��z�z��a�?�-r[����;����O]�2�h�J����} ����3�Z�7��j�F,�C�E�m�>���b��s��#�p��4j�M����&���m���L� ���ֈ���6��3��[@�=Ƕ���p!#����/Y����)��Nُ�v4�'����9K�������c_��G#��/LlQ�JUZ|Όy8�����"$�(>�a��w�İ���>.(�Z��O�J�g2d������Q�dU%(Y�ND�X�PK���������Q�E����*��乭��;��c6W��攋�N����@o��Ku�MJ�ƔtE=W��Uѐ�Dit��0�2�Vw!l!U�6Kڶ����5��&�9���A�%}���A�'��xsmƔuԌ��G.9e7 1�A��ac!Ý����0C����4@Fl}��@�}o� \c�Bc��Lf'�!#��:�94��`;a��߭ھ�0*�H��t�gT�nб2�"_#�B�;bn��w03P���d�Q��e��#y���JK�AU=�3���'�� �(����SI9���
%�aS�x��H�ЂQM�����p",�D�<s�}o9Q��:Q��e��"�S�F}���}�8��M.��~n����T^m��R��@���C?�£��E�E��VhQo����¡&���Q�5�w�mV^5�%G���?�?'�q2>p"7��Ē�;�";z� �i�[
_~���%/���m��]�^[G��VZ��@	���Un�N|��� knΨ&8�ݢ�t� <X�ӎF���E��=�F�yB����Ұ7���X�7�G�flZ.����8Q|���9z[;A (NH?#rֽr��� L�4��،^�\��iS1U�¤a��EQ6��&1���4Z���l{����;��"���J�s���e�,���GKC=���ӷP��!�'ς4��9jˑz��?Aֶ����y�����Դ�c+ь�(�8���޾�t�U��������܆�g>���ę����k$v�QW����/?�m�����A�j�-��<�1%S�5Qy��J1����6�(��6��m�B|d%]:�alA���;����4�D;�Xɨ�K��|9�s��'/��&Hx7g� �21�1�
s��9`�A
ԡ`p�'�Ȅxi,���M�ry��e8P �v91Q�����!����DI����y���as��@@�!��� �e��hǾ��@��U�-�+�
�+�tu�f!�A�	�V�$.cYA�EԊ�N+>��tA@�񧎥���xL�Թ�:��*�È��E������/4�1~8�?�X��$��8h���:"vu)�3�6����UJ$�Rq;�2ŪJ�Ä�\=rZ�ѫ�kL�(��l��?���!e+��n>`�!��_���L�	hM|�fS����I��5�T���s��B���q�CN3�ȡ�Ұ��]#��F���g� S")�
\�kH2Xn���ٷ�=䌮{���B�v��Y���0>��-�e�n����2�,��*`�r�P&%g0�Z�G�E6�&����Y�+��!G�hg�n���Ƚ�E[E�b(�6�.Q�[��Vݟ���{�����DU�H�לּulm`��Z��DJW�Ir'$�r��O��lx+\�]eC�
�"��(m�>�c�<i .��ݥ��6�񥐐�'���{�5F�d��r,������V?+Lo
��D&����e�`*��$�:6�c^R�m�&�MY����	�����[�)�y�5㯂�i�F$�\J������K�hl���bv��v'ˆ�/�^JSة�Q���5./���n�1ǐ��@�0���h�RŀB$h��?g��	X�D\6�"��c���ݠ�z���A��;��\B�չZu.2��F��?�g"�=}�*L�-Z\Z0���%��;��_���I-Zr���P���su� �z��%˖*�,�D����u�����Iu�$����b��c
�s�3����*,	P&4�z��횏r絅�.~���}��w�/�������H��a+ƛ�t�B�����HN=��:��5���N���H��\�Ϣ��8%lBAr'R�FTO�9�/n�h(p��	����/�O�/	��g��q�TL��tQ ��{on}��0s�����RG�4<��A� �P��`䢨�X�?�_�N?���zN��{�<���'�C֟^@�W8R�/{�զ� ����/��J�rA��>pc/8�cWd�!!������N�p}�����EȄ¤����//P?��1jͥ7e,�yS7��+����R��R_�d��\���oۤ���c3�l�${�
��1���v-�}��⫿F�
�c�@Ք�]��ɳ��b����.l�vp�QT�|Q~��������yڍ^�F��a�$�����׍i�
��\����.}�H�f$<,J0���y��΄�JE�?)V�ȇu����f"�����P�Gb��g����`��3��D�Lf{/S��Z�U	�����SV����n�����������C�R�������e�D�]
Tv���sv����f%�7C�2��=8�у�J�hl��-�����+t��X�!��w"�Bw!�cF�a#���Z���v���t�k�N�x��*lc-�b�HpqS�'��"�]>�������(�W�}��S۳|�����;Y_�u}B�]�j��\0 "N���U�����/m�=[;���M@��z��Vf��?�+n��*��{�^��G���א�dKKY�Ou�kn����<P��d{�i2w1�!�R���~���t��:k־~�ð�����o��K�d$:0���D#���	D������´����o����[�8`w?\10š2�~�D@�0�͝0�)l���"t�>����U�d������e�W��^+�3T6�s9��eH�p4IK��R����������NQ��. ���u��J�q��'�d=H��K�c��q[gg��K�߃`O��`���e���߃z��x	��,��麓!��V��Miwf�jP@��Q�Ȑt�zr��h�'v�x�.�U�A#Ωa���|�}[G��Zq� ��.J���a��D�U�
������pxy�'�\�6�v	�J�a8ӵ�G[�Ѧo�>o��s�9��5m�����ͦr""��1�"�~�v���^�z-J�2gy[�xm�F$n�щY�,�y��-�N�o�X����ΦaF�B�ZuI��a�툌XNo�J�*jtDo��&��w��9_�Z�5���j�ԐE)���ɦ��Tj�ӲѤ�C��U�Q���ظ<��~1^���fu�U��n�Q-~�j���l�+[�#:������Ƙ}�}�tK�����\"�8'�)���p�>_.��ś�*�Ru���"E�u�׻�lqMZ����ϭʝ���qN/�璒
ynE: R�j�Yd*�l+FdG��mŹ�yS�<���ƃ����>*���'O2�-��D�9���3�&&��6�]�P(�n��J��82�s���?x�H��FQ��[��a������a�G�K���X�잂$|��it��V��1����8�kc�� 	AI�iWW�(����E�̦��P���B��hO�qݝ=�{��}�"+�d�i?9������T��]qg����[�U���?��c�tb���R%���n�h@�`ԍ���y��풵��*�-4��u(z��z$��Ma'�C���ut���p��A�K����^������=�L_L�|�H�KO��\\�O�!(���B٩�'�s�ב� tsY�y��X��+I��V,��L�ݢ�H���=!|*�J�͝���c}��^�9�@�Y��I|3�֝l)��F^�+kwwRN�U�n����ي��^�����R�����EI��1m�G�j�*_�`ĵ���mJ�tӠ_e��'3��f:"��iʶ���p?��
�y��i�j.���_�z�>u�k%�è���n±��8E�V>+0p����TK�}1��Yq�hԹu��i�5��q� Q�y��91��]��ב� �SU�Ao�+z����M�ݢ��c���_W�<I�5>��B�*)`� �b
��b�4Z�Gm�t��M�."����8zǑT�(O�hi>A�"�v�=�/��f��½x�������Ϩ7�/��AQ�ڼ�Y�<�^�l���.n�-�}nog�cI0T4�C��TY�	�UE�+�6��G�m6�[��8������e�8<���hvP�Zآ�#��Pd�mʬWJO�s�r|�i��9�F�i��Ɓi�|��1��ʮÖt�o����Y����Dj�ɭ5����[OPf���F�Qy��N0:[P�m0`� x�w^���
�%^�����o7������T��!��`�%�=o�Du��s�������)���'�mcc��N#i0����ŭ�\�f6��튧��vXad����	����6������S"Z�Ġ��W���
�Z$�5���iH�D�Q**%���H��=��|k��2I��7_W[uI���n5O���]jݭ���H�c�O���j�/Ͳհ����7�QG��ʄ$@�ۚަ��
gњ�qB^��ڙ�4�!�q �Οth��JX��$��M�n&��۴3�X2��󉓠���[�i@:��=i�l�KS.��A��$}+e;z8���0��|<��\����5�\y�Ϸh��.���kr�=Ҵ<#@\ܪ%���p��׉��л� yU��z��n��h�V݇l����8R-VC붍�I7>=�-��Q��6S�Po�֛�S�K����+ihpZ�����G����Pf��b�~�N��×�xƕh��=`��gg������+�q�k�#�\�
^�{h)1	3��l�v\��Qv#�V�:O��!W���A,���^�2�N��2���ʗ ��8D.�k!�oDƿ��8su$��P��;;s#�kL�Qx�ɘI�G1�(�P����S����p�c��CL&=�3R�'(ޜ�Np�����/�w.��PC��j��BA���G�Qh2�� Ӯ�sa�k��Ne�ĊT�3Aے����;�u ^�J��ʉ�y�ʓ3)~�_m�2B��vj8^�蜂;7×0a�L��c�2� ���];�n_W�0�K��[�ͰL1WiJ�C�cut]����$�y:y�k��!��L%V,z�-���\@����#�mM��_n~51T|�s��e��<�Q-�[1arv�?���6���g,�b�TbS=������6���:��Ƈn��F�������v����.'�����_�ç��ʠ� �뻄z��%�g�ޙ~�ݹ�R���u��!g�yw�u�9��l�=�'�n �l ܼ1�=꬞ã��0�W�)��`��c�@e��� 
��ETLWܻz-	(jd�Ѣ���,�j����0[��]�:W��_��hӐ���4��K�)�L�S��"�6�*`����4Q��j���(r��L�a]F�?�Z��Y�:�qƏ����qV����k�ΟBw����K����j���X���E��Z�.���gN�ӣ���S����2�uR�T�_�S�~�4݌R�y|���	��!��������]�-l3+�x�se�f��V��gӸ˸�����U �%�r�����Ƕ�����l�'���yP&���br$s��>\6��z�����*=�qc@q�&�\R6�ի��$�x7jG֢���{��-�ߐW������&��^�|���&a4���NC����o㝇��Eq��ASc�v�ǖ����}�r�k(�"S���,����h��dC]��f�D�_��� ������^������cֶ���P �@5�N1�Q��_�[�7ڶ@iR'��ʪ��zIu�ѓ����H`]��g��~��N�uh��f'�q!�y?�5��+�L]�	��iˇ�Z.9�T_U��ѐ��OFX��|h�x���?d��Oo؟��<��	�����>�ݳ������D�\��Qv	�Ά%l���|�/�Y_�>��jDRJ�2QDG�%�n��l����p�xX��G,�},n�w��Ü�����K�:D�㕣�#��s��	�*�RJ�5����~_�ٟ]��w���<�Đt/�*�^ �'��U�Ի�~�6z�мq%�Zd�v�M���m��f������v$�	"� �3�C��%#ܪ}!�(��Om�)�K}���\�*�5�����d�g���I](�y�͇V�\5�#�1#(��4�32 YY�JN4�o���Y8ԋ\;;�:W��XB�ʓ��v+{�O�(�za�?���8�4æ�oXG�H�8�Q�#8�#���1�6W�.������	a��]��¥bH�Y�*b�jY����$���qZ7����n9�>��D���&�[��//����U2ɴĴQB����Gӊ A�U���@Ƞ۾:aý�k/yY���m�����yj]�<��?TFm�)!۝,j�����d$�
L�j�y��3O�ir��\U���F�n�ff�!r�F�M��&ޝz"�W�<��oF���K�{d�=���1?0���/���(l�pu�.Z�4��jFیr�o���BN;����I�uN�}
:V���!��V��#��HSU���X[�����U��@/��l76�~2?�c�AzF��s��"�q0����؃{\�}��Cy<,f���8G�A9��l�8Α��qGPV	�X������fQ%B�NZ��Pp�H��8�0��aE�Y�p8]�"�_�yS{����%�?�׸�Րj��P[4�6��pB��b<YɆ�M�wn��>�3��� ��_6s��#�w�l�<�2N�L��BK�	����\�8}�f@KV��Wd������!/ j��M셶��$KD&�*��}�(�Ë��}�w�!G��Y���*i���f0��U��	�2R�b�a�Y�.��@CuX�(m�*����ŵ4�0;oJ�h�-.���\��Tp�m��9�T���cO�s���7 D�Yl�GK�5�Y��{�PO*e����q�_x=�ѯQ�K���@��2����CFxw��n�����h��	�IE��Z����[9eu#$kD�#ulZ��?���ב��"����H�-J�KRpw�a2����=B�v�����_<I���U1n�D�-�D4��kǿ
R�z���.x����Ͷ}�@NCQ���h��cm�U!Y���?�����}�V9`�x�+n�}��qw{�G^� �uMn��;�o�gs�p.��aЭ{=]^�m������G)�Q�t�drǩ4�`\�"~�����g'"���r��E����K�S�tKX_���/��3E$J��Z�Ho��D��H�ב�ј���*���ctW1G]��ƍS���B�M��QW�R�zQ�FUs�|�G���Z8aI�=�H�>�s��Z3��<B�yȯT�}�P�6H��"ߥ���2>���5a�Q�p�2)v�@l�YL��e�x=�.��縟�����#�11��v�T�Ty���xRo+4�v� `�5�}�G�d�u��Pi�,�`u�0���&�*u�����ɴA,X݆E4z��O�U{����n�h�Q"�Կ��A�FbtL��R���m�O�-V5��C����&/x	d�MFx�m�x��=��t��*���<m��|H�c��֍d�}�dD5�P��w� ���l0BI.(�
��}�a���8#б�A�Fc�xn��D�ɬ��FBmvg^e���E�"�$��~防���	'�B���ՐX��7�s�ɬ6I�]����Sc���u�,��@�\��'`��C��oB�f�jQ"�F�j�ڧ䗱ǵޖ� Z�;3���S�}	��c�u^�)E��μ�Cs�d����Ǳ$CJ�35�qZm�� F�e���1��@�T"�h+�;P�l�,jh�v�DAk^,7�+������E\=R�c���3��}�-<L����ű���_�q�!��0���N���4��Z-`�2���X����T���DY�0��rn��:�i!�>M�ɈeS�N
���67= Ug��)з�';���ϐ�'����yc�ۤ��ׇ��E����﬏���{��f�$�Hx���+Q#F��4��~q���~����YA��+*�(��䁺6i_H�׭�ud�� �P��y*)s}�{�Nx�,N ���m��lY���d��K<5꒸��m�F8�۟8
��/�u�,�P�d��0��x-�g�z��~�I�8��߽}�[v�<חcc&�S|�����lE�VH`�;K���;�s~H��Ӈ�đ%���R� ���1��m�މ�H�t�Gc�|Q�%N�G�C�k-m��y�L�4�Ԇ}�¯�'<�h��w/�d��7o�Ū��}Yc��_kvGI��p�S���+�w	�?�K���[6n�ں� E�o�^F��*�!#�rЁ����V���	�T˥I���$�=�m��`�E��l$R甪��Pʹ3qȴ�ƒ�ڔi0�S/�Ӭ~�0����ϗ��=O�$�v��2�O8U��G�r^ŝ�9q%�w�Tض��3IBݛX	*�ʘFwmӎ��
�������rՊ�deM�=�j��o�",��c�%�����U�BqX�x�N�ǣm��:l���7��Ks��s�X������X�����'s��2�Ҭ/�"����?�7ф��FE��$�}�aܤ45�EJ���iܬv���F&o�ڵ���F|��N��2���o�	�����ԝK�a�*ca���f0����yɠ�#�v��}���P���Z׶ĳ�9����J�q�[��Q~,�iC�f�E�7"�,��;(�g�e6�
�J�?��$��c�o~���m�N�E\ہ�KY��$�C��ibZy�3v�]%��%If���9���� ����J��#�"���݅1`�����xt����P���5>;������P=D��b�FcJ�����@�SO.��o�&�<���E��^I���D�QJ�t���l������:qP`ԝU*�U��c�L;���<���<9�Ιd}���D��o4(S_���[���`eXf��9����amt]��{����Kqw��P\�k�'hqw.��ݝ�R�����_�������d�\����^�,pCD=���˸�C�[�&���r˾��)�1�6U޻�}�G���\;�=���r��Gݔ�L2��������reo$!�fW�Ǣ-/���ũ�κܽ�2tHsg���eo�7p�����O6]V�ifT|a{�gCIر����jp��
����C�˔��5;�!�ٱ(0N%{���+X��遲�b�˅�h�F�V<��NaFv�mZ&�,��^�Wqw-S��t�_=1���}�
�0A�P7��{�Ș��5^C22�}`(�_KX�)����������+y�,6���>����u��==�'J)�ӬTE� �8u�!-����ӥ[�/�7eT�},��?3щZ���{��[�dj���Q��)	cpj�5��I�j�VG�ѳ��[��k��K���	[U�M�� Y|�J��z�����v[��6@GB1Yk8�r&"�/�g/����$�����F~���SJ88� Kq|���P���A�𵸊|\���hL��.�Y���ٴ��	R�T$��<Gh���Pm���!�|R�u�O$��:�d'������k�L�,\����O>P�6<���Xl~F��?���QD*��&^�*
5�eE�s����a%|�֚l�a�D-�aߢ�"�i%�F��a�+j�tB�I�#�~��;�垣�k��'����<p|�Ӌ���?�Z�-Tq�e��K�(3m��k�YK� �mI/$�H��t+�+�')d��	����k�(��L-�e��}dk����o�����e�Oy�lB{B���a$g	i%�V`�؃��Ȳ�$�BS�T�f?h�]����ɞ����%?`EY���Jd��$���G�L�ѧR�BBĶ�G�������逌>����$C�y���d<�}�
:����.���[��	+��m}?[�_֑Pc����C0濛��I�oh���JXd��еDF"g��'(Ӱ}-Z�B�R(QGƌ��V��?تf�6�C�0p��W�ڳ�8h���7��YVg�P՜ÿ#~ic�Y7��[m�����ATݹv2�Ke��{�(�js�A�N|M���]5B*��Ŋg���U(�»"�8g����K���p-҇��,���ܩ����5[���)��К/�c�OP0wTg�Nm4gz��~&��K�Y���|Q���]�;�C&㉘4B*��Vmbmc�3�O��@�6�٩3s5U���ix �ݭ��0�DCw���� ��Wbz�Ø ��:�&�����I�uk}LS�#n`��e|
�7B�m�'���p��'�W����f��+�����>�-[%�ۺ����{�v��ǭw�6{ŏ��D���'x}�㘕�N���K���;͚��r02È;���W����\?F�=�[��	��}�C?��BlZ:�*o��4b�wѹ=��pN#w�t�Vϼ��j>�a��|��>E���l���T�!&;��o]��ɥ//�m>@�=	�\�R:�n2L�����aB���X���մ���[ƶ&Q�۽�a��q��p�j��	��,nn���n�tZ���?��P��Ϙ++ͭ^��Eb�c���+u]/F��+����-�!RSG��6j����;����F=N�/^�N��б���x��5�%��k#+ط�U����XF�X�G�|��r�*����j�A�`<��>!}B�b9_�r`t���}�p��b�=K^Z�����ԡ��/J�Ɍ*�a����nq2�����[�P��������c9�)L~;E���}�N噯[��4�D=������<Y�f���z���
WD��̟�q�[f�ٳ,:t��+���Y��p�2��z
k�<�ٗcE��#��\[�N��W����g��٣U�j]V������Ґ	{7&��+L@*:��^G$���y�"cy�G��X�
ƭ�V�cn:���!4����V7^�3�����N���,ƔQ۪�D9~?!�I���x~�����]}�!�v�E�Yi�����C�t���_i��vU��^����Ԍ>u?І������e�ZQ���+����|��J�%!ٌE��p�����zD�!0'�׷��o��c�rI�$'��b�⬫.h���/��iɟ�8Rt�����?��2��l��������*�HO]t_�(��.K� �9�r�'���?��Yfz�R`���.0��m_��_�&��{U`Y��K���p���@��i{xY��mq��ڈ�+�Ȇ#�R���j�"໛���K8�����Ա�$N�����6�%C`��t+4���D�\ع�PY�y����"�8N�1HXe��q�E�xV`E~sw�e�cӿ�睨�W�`/|���%�|�����}:+W��(�nY��{��*�^���F��
�c�W!&/!䗓\Ěc���߫�����@��>�`6*QP�a������]f�|$�T���d�~۱�lM��`�"�_k#�%�A	M���T\Q�N�l�����~;�q�����f�$wt�KQ �<h6__���>�w^=ߵ�ˆ�Q|�Ʀ�"A;Lҭ!����,[���!Ya�+p�������]��D)J?�5��j�t�T�=��Z�{�Q��#�dfûϨEs������չ��(�:�	�~W��=`�d����Ժ�û��Le��Qo���WJ��\ ��<�@t�7E^'%o��H� ��={�����w<�Pf���Q�Q�V�+����w7��\�� ül��N�3�W�	6Ӡ}Pq�%�DE��J �,t��F�XL3OY� �Ҷ�GiUrֲf=��۷���f�>Qw:�$�P�h���\&��k�a�j1�k>�^��ف6���d�����C٦JF58Nz�U�	����oQS�ߋ���T$�zU�KZ�;K�*oW��$JEw�N'�1~җ:�}���	?�-%��HgfF\tO4.�֝SQ 	[8��b��9�y���b�FGU��[�6�e���&ޕ���ACν�<�͈�,܋��E����w���[Z-[��y;��RX�T)]?.�*�e]����|e���Ã,��%�2�<Q�11��ZZZ��hڬ��uݐ����x���}����y~����>�(�`���K�.E�@����t�儢L;���Լ�j�?�L�;���(��ZoT�LG�3q#�b\��Q�[W�����ֳq�!�Д��eB�f3�G���0'0㎮NU�	�N|o����ѩZj�˱2}R�=b�A̲뛇���;�4��*!�C��{h�����mcES�Q��U���w�M�����>�r9a5��Fڸ�w.�:��,�E��*�z���%9��.�� �Y9�>(�1ۻ�*����}����kߡ�p�x�_��y<�� �
-ܮ�{a�EAo��oSތ(F=N�����^s��Y��*i\>�a�L�L'�w{�<闌��$���ܦ�S_�>��R	���AY����Ùk�����CQӘ�f��m�����0���*L��,h2�4�� i,��FV䰮���_����Ú _k�����E�IzLq��5�E᧣[O��ܝ� ��O���H���5���We=��#��.d�[0��A~og�o�Xd�oA]Rr��������N/͘�ک����$+�\���t.Q���ȜB�K�K��(Pc�bq`�?�Row�ѩ◀Pm�3)� �q.f!<�{z@Gt����A���^h��Nl
G�+΁�|��!-7�+ϻ '�I?.�"�
ܱ�:D\��ց[I����*N����о�q�z6,���h�n/�����Z�M��&<��M�� ���b��Q��o�K���wK��f�uj�գ�1�����ҷ(#�^�2��&c��E���&i�v���Qַ��lh�RŪ�P
U���ƛ�b�G9ݼbT��{k�M�#�IT���t>&5i��xJ^�����I�l�[�}�(=��Ư�gh6X�"&!���jǸ��wN�|�b��/\�pZ/�09�}��& z��6�3������>��}k-�f�s��H����^e���\ɤU�K��2@�ěݓ��bo�iｈe�߰�˝>w0gnӒ*��"J-<X(��H��1���=u��Rb���٪�����ה�V �6���>4\vz���5�^Û���W�RBՌF�3��O�ۥ�f�emC2죁Y�AuD�쳀�)tbO��>�G� 㤢�Ɏy_��A����<�E��GjϞ�2�����
�M
�|���,�s"��(V#&j8L�������y�!U�\�ZV��߆��"s��U�>"��W�o�3qy��}&���B�l]�1��;�V�!�h�d��J��l��8h���j!���;a�����g�o���;��U�7�%QB�W�߇n�R%)䄵��
�{��ѢR6e<�~Q�O�C/	곖4�w{qq��ڥ@"sJ��/VL?;�n��)�d$��]��9�>�-�!+�˩����Ho�A;>��z�)�?�̴*�Ԟb�a&t;��5�Hk�7��7:~��9X!٠�5p�gd����|M���z�s����}k�>���0�jm[�&�vo�q���d|�Sq�����V-ps5^�����eYZ���ҢY�^XUX��U��O�$v����)��D֌%���M�a�?���I_W�'�S���]�~��#e�o�,�.Ք}�j���}�bd��YShll!=��3�Ąp�)ϝ�!wy�c��",A��1eq���ɠ	�R$��]԰�U>ѭ���ħ
�\�N��I��+�O�c�5aa>��с!W�!=�gPwbyf�~HR-���X�0/�?��"Q������9+���6�?]�Y�۠z�z�5d+�$���CW\#7�f��e4~Xe�����/'ܳ*+� vqQ0�=��bm����-N���m�Tg�xfK7fy�[��2��랊
�z��+րlSǅ��ۈR,�Ǐ��l�Օj�B��c���a�&t��20C:�Z.ͧ�HYVz�U|��᥃/��4�hL�����m���]{,9��>� �Y!��0α�ʺ��F��!�w)aO%�+vX9I�p��ߣ�9B���f�],��O��3C�J'�i8�*�o5��>�|�lH�+i�J��r�P'��î歹�!8�Ɣy.�A���i�|�7��kOƨ�mc'-��.
4���wO��8$��κ�SТ��/��Kg+�:���9�)�.C�|Q�%�mY��<�T�sV��G�h���7����y�F�A��ہo;�R�(U�O�ҙ����<��"
L��, j������VĴ��Ԉ|\(e�҇�x��ǡi%ޠa����b7E�$���h�E�S_gfߎ�P�%j��r�	2w�7nZ�ȶʛ��p�"
�.~��Q��ٵ�r���I��d�k��/8���S��JDk��P�K�0���J�kn��f�p��������s~�>V�H)������$�6#9����A���d"��S[�W"�!p�pL���̽��6�-�u���p����D�K��p��)vf�d��.�$ێo4,~���`MK�����-� \8nԩ/����@�o��w�]]���.S'LzP���lB
��� �z�5GLc��n=��)�(��Oj���Z��LӤ�oaXsa.�u�Ȃ<,���������)��gN�dj�����̯��?}�:D���ٌ�:L;��z�KA����e�-=��Y�Ǩ�ƹ�W|+$k[�$��/�_իoRݵH�y:�]ͤ�4OեWٶ�}a�v�+�AGӉ�Aῼ�D
*&���aL�J[�g	l��+Az����R��Z��"S�#���ݒ7|��p%�f0]�|���^���p<�xۛb�Y����W
c;������H�ecG���b����벏|Sk|n�ƈ���� Py���K�e+Bm��9�N�*3��k�6;r��J�h��[��4�f�6��?5�0�e����?��K��� E%�<4��3*?�`�Be�e��y���D��\����)�p��;�:1ӿc9kU��q�a�3́B��0�_ׅk�C�$�۷�c���)'s@��գ�g__�o>v����	�����4�c����[vv�pM�S����&FK%SG��+	��4=���g����-u�����3Q�-�/���D�)ّZ������J�O�Б��d�9�7m�>����%�h���J�Z;�r��s��l�¡4R03�7C~��Y`��"W:����}BWgL��V!Y�����QO`�_p���L?����e��d�h�
��Ѥ�7P����1�=<J
Hst&؛�a�gw��@��mWQ�5�������Ä�qYH�{���;�(����� S�c��9w�,� #�
��g���׌m֐x��`��>rs��KQF��|����o�#�o.�{�����;&v�㟯�Fk?b�XE���p���Z*�S��r��v��ޔ{uʆN���xD�d���!�Ӣ&���A�0L��i�B����Ӆ٦H'_�j���V�@iLkWU�͆;>?�ܛ�ȶ5Z��C���[]B���B}���Tg���%�[8\���X��emI�<����=nea���{�LL��fg��s�Z`m!H�����M�H�	L]L���Ȓ�Ǯ�H(N�+���J/��'�^쫌��٠O\��3Qi�v`���t�$M�9ձ��Kȧ����LWL�Ē�M���5HW��#j��BؠI�|���*5����C�$w�,bM�a)��̧��"�)��$g�ɛ��g~b��s�Q�ʧ��%�u{T
Y�q���x����e!���@������j�����2ռ��}ύ;�>g0���~_	�^kq gEb��H�`�)�������O!G�A��h^s����ٽ$���%�'l�����)M0�	Gx���ա4��,`U����p��
A7ez֕�z܃���3�pn�kS1z>,Tq[}ў�s�u�*�����a�B��'���=-�E��"��xM>�����vs={��"ڏ"�Q{�����|ˮ>rj���o�⿵ wڊ�9uZg��{w�OK�_��'xg�X�����������s��b�9��t�Ac�w�gv���xV_H��߶8s��ɼ8�ų����
�_��l�h��M9��M˲ct��7u�[y�|�V��.K�'�S��xv���0��C��D�i����;7<T4b�-����5 hf�T�ѫ�c��Y=�ŹVXQū�w�m��mF�&kJ��w���V^�gמ�t���5�F��M�L�*�����u9�zn��~��wdnZ$$B� 9��E9��N	�.Zpή�P�O�t�?(�"O�CC~%Մ����ߋ;"��>p�4>�yO���PY��0�Ƚ��A)��`�CT4'$���h��p4�S�y]�`���U��2m�N}�o<��T��b�,-�O峱��'iJ�L�H��gt���`�&�~��[��Ζ)DL�:�Z��=�O5�lV�<6��6܄���I,3�3���l*b��x9괛7_*�lR{��*���]�B���d�!+� q�yYdJ�̹	���1�^����k��pTcy9����8��1��E;��u�|.��+��9ֽ�*rD|�0�4 �#�l#�F��ɭ߰���u�f�zq�u��Gf���I
<�(�EU�>#������!+V Z)(�������ZKb>�k�j�;�eLqͳj�RjLnj��2��4}�İ�h���� ����	�EPeDȸ9�_ B+;j-5����T��8�i�3��Қ�l�S
{m�U@ٓ`jys��D*�=�/�V�o���q�E3�J�r'
�ukL����
�`?�O��)���wE�Ya�	��~�
�<<���@d�kɱ��[��Ls�0&��ٗ��K�|/f!wGwO�����qMXBG��U�i���}E��������ߚt��t��M̃d�L�_�%H�	������J�m����Gi�'�'�C�J�,�u���˗�Â�z�o�P{�5�J���������x��Һ��x�-� %MO'� e���C�Ā'>��[�����(��ߋ��u�٠�ɮ��������Ƿ�c&�0�<7M4<�Z�)�� �C�AtǱ�%�O88/���dAM�V �Br�OTu�N����yj�Bp�G���Y�'�G�*
��g��������΍���W����@��+o�KJ֯n��bL��Ǚ[Ά��|d����R�T=�F|B0n��.	ְ�#42~�Y@�%ヅ��+�c�[�o�9�I�5PA�$��*��9�7��T���n6�?4���-%0�>�|�(�hP2c���L���DiQ�-�P�5�`V�)�����'�ph�ɲ�o7�T��'����xf� 8O8�f�#�U�ئ͇��b���C7?��b/����7�@��]I�P39�D48��(Ö3^����6�A4�Mp����J�/��܁'KK�7L'��lb{�/�0��_�i�r�͵��n͟�q��`ڟ% E���Ru#��}u��YW��ˤ�l���Ѝ��0VD�x��+�c�'�'�9�0٤{��PX��g��� M�~�B5b(�)�W¨
��՝��
L�h��T37f���Ү	>���M�G�T�H��E�������hъ4���d?V�����jM*/i1r��I�(��[��TD^��c�}��ѫ���e�(WڐO� ����v�G�0r�v�\��ь
�ڐ�l�_��:RZ���g���|A���Wh��'kc��a\)����N�{�:�>F��fT�!��!��h��f��*���|P��*8��[p(9bp�ʀ�X���v'�=� Z��D)�̃R0:�X�)��9��y���j!W1;�" Ȗ?�n�^��o�gt�N=���X��q=rKB��l���G"p�����Pᡨ�I�&l$�@�	�����v�G%���o�꟢�khU�?>����3�maH����d[����!a��]�_ND:>�܇�v�=�_d�Ic�E;�` ���$�r�*�	{��9�u���sE�aĒ)ؚ,���[�w�A{E_L�����+�tfk���X?'�bHZ��bgL({���=Y�b�7Y!�ǔ~�Ճv�&)a��ǝ��+��AD�D5�33��/�;@39���R6�ݷ�Q&n[#$�^���=�L�l�t-�K�m-��_�G�Q��6q�q'XK,��=9�(2�(Kb�&1��oˬ���`�r|�Fg���=OCV㌽ ���G /����'¿���H�s���&�b���;]�'֝�s|#$]���lfy_�����)�\�'`cwy#�D��h�u+.|��1��&�~"�T�Eg(egF��5�·�`dA����k�i\��������#��j2��+dxmp	�S�j����"��2�y5a"���珊� ��ђ2Pj�I�F�Ա�wz{h39��D�ͤb΢Jнz��g����)��3�]h����bk�����O����#�����x�	1�3,���{�xʮ1�����AF"�Ieƣ��Z��v��NB��mNY�c��/��I���˔M�Q�Y�Qp�4���ǳy'�d�M�O�w�v��� �R�}��9av3;�)3�W+�ϫu�zl;�;ŒR�L9U^<��k#`)�?����m3�����u��č���:) BX����粁�y���U����m�)��і&�@ �矟�bg�]���=��L�~ް��+Ej��0��`�1�$F��,�8�\Vy�^N��A�1�z�R®Jmj�t�U����p�����Ċ[�	��v����&�澨T>���7��J�*�8J��x<W=~���ϑ���3�O;���o"�"c��t(���!���i��,��takJ;��ݫ77����ن��H��B4�z������b�ħ�D���uhT��� �ZH���ж�΍)sD�q6����h��l�9��8��u?���2��|`�����2T���^�}o�n7Ş�5w����L�Tx��CQp=��|�p#�:C�^��/���L�qB���7xѪӥ�z��N�#�5�3�+�=�����+Y��mT�������	���]~���*n�9�Æ���^�SO�qv&`:#_�Ba�NWtz+M�Fb<��ŠyM���~�n�I��݁*�z���B���f@(O?��JM�[�^Z�@�[�`hCz�u�׮��i�����ӋI�U}�_�h��e6j.�t�	e�.Ϯ{�=�!� p���]��9�hκ��]
���e���2� �Uw��*n4�ݵ�A��<��[_��f�! >��閷�/cW4?*$�x�`[��Tʾ�N�G36U{��fܠ�J=�?jAL�$7��P!���k�T��.�y��l}]�gܑ(H�#�&JԘK�B��vf5����_hC�M�k�d/ڎ���MF}�6[���.^��t_�G3��L��(M��x��O���ɻ,!۟�W�+��D��$�s�����C;��Cu)5�h(��}e��Gݩ@Ą�#�!�b$��$��t���	:>�b�e2���vx�����%�%8"�@qrC����먼n^fw`QV��_"��?g�1�'^��s�l�S*�[��-Oԃ��l䛄��-*�ѽ0���淊��������2{<s���4��"�d�g��aob���P�F��Ķc6&��Q�!���D�����2~d-�H>�+�B+����L|b�(4
��%���	s����R0�W߹z�*�O����X��-��0?nR+&O}��Q��t��^�>E��5��t��+����n��s�κ(���/��#���|����6�$y�q���Oe�Q%u,� ���V�R-{Vu�E��ѭ'Y�.��;ѿu�J#��5̋���aᴛ�p��Jd�3�� v����FU�<G^fd�߇�}!${�%YԬH�Mu}��o9�����9��/E�=�=�(�����x����Ǐr�?g��6��x�n�S ��c�b���v�h�~>_���f���v�%���+�-�˯y��Z�J��5T-ĒѨM���	^��	���cujD����Z_8ʘ�b�ҁ��^JƧTF�^MJe�(�YjW/z0"ӽ�d��*���f�{��>�Ҥ���I���M��V�t�fbN����g�ML�>��,�&2�2x/i. �~(�zК�_̸61��]��4���̉jd	4�����# ��r�Ntj&����+��Đ�?�%�NF:�5ҡ��"rw�i�m�A��J�`Vvb�r2�+�/ )�"��KX��{���)�e��ԡ�����k5uq��V�`j��%��GD�_�W�
p/�[�I9�1�����$�+���(l��q	�H;��˾m���^f�g�2�������'ʰ�{oQ�?L��$>2s�z$�W�qL�`즗�4}�[�`d�cH�M��fL��LW� ���v�[P����JI�UB����'�`���~�
 �m��G�NT�z���z�չ����
*�(�bk��}U��6#�����V���㹸�\��:r#ӟh�tx�8Wi~� �Ô���;.�)�{��iPׄ5gK�����3�5�A�L&�=��q4ǩZ�{�u_!G�:�o͓k=���c��炽T��/�V��#�kQIu=J�1�rs�ί�3������NJk��i��j����V+�E}��C�L��E����R���lI���8]K�+��Z�nɋ~��0t��l�e`k�G����GORZK�&@c�A���ߣ\��-ЕR��'�2�yH���]�	h����>3�a8�L�K����ҿ�ME�+�Y��Z��f��4�I���I�ۓ���lq	�g�G���j#��T��HJ��ۀsB��J�K�����C+Nd�Y$B��_c�GizG-rV���E?}��U�hX�BH �5�hT/(�r�B��)ԇ��^4S�5i����EuEz���p��ĥ��Eha�C�*;���q�*mNP6=���������Z]I\�9����q����R��7�V�7t�u>`;�efrD�q^F�|�����#TkT=(�z= ��h����/�t��X�z�}$RTxMG���{8�,ou�����pT�h�#˖�@�W��h�=�C#�����]@��H�C��^>m���i�w|�vj���1���0�.3�K0k_%!#k�+���:��g��g*X���/���,�:�i��xL���5��J��O���L&�s��'#Y=��3'/�pTݙ�|&q`�3&+<r� �
5�H"�-�K��A�L��j�s��r:�PŽ��0+$<�ʙS���W����'���]���+���{m:	�f/�3��&g`,�n)��$��5�IP0쎹CP�Fu�&��Dt��u��]>@�}�*�4� ��i׻���������x��3����C�'=��
�U�ֽ�U�z^�5�ϥu�Tk�d����:/��9G`w��0�N�E���u���&ə.�dO�J�)���QA��d򑎪�H;���~vyfu��H�\5��ðP�BҚ�c���Y<j��<����
�b�V�u�V�3hf]1I�+vT��ve�V�x`�hk�/iT%�y4_�𝿵������M�6R�v��2��u��m����;�*�h=ܯ*�0qs�v�����m��j�2c6{.����(څx�I'Z�5Uf���ax�5UNT��1�B���?;���o\�n�{��"�|��������Z�c���	߷*m!d��@t�ᣗ|�{��mTP��)'z~��`:��bޯJ�Nw=`rQ	m�����t�B���w��v�)�-�[p��~�b�|$D��GVU�������zn��Z�&��毝��?��d��H�Y�bE�R�!��k� !6ǵz�>k�������R��YڧG��d%O2�s����42M
�2'=�?nߣ�0��ƙ����������Hޖn`*�^��_���m'���N�.��Q�s������ܟ�_7�7�K��A$ŷ�c΀��ň-0t^�u��nѕ퉞vK��w�"�8��@�R)V�:�=�X��x�m(��O��� �{��s����4���5<L@"m_n�M꩜ִ��'5�l��<�'��`\}��0ƀ�^���]Dz���Y�.$7Pvܔ��hm~in���e5��AM��'v�����l�a�.P�a�g���և��{�l,���@��﬚�>�Yϟ͖�U	3ip��1����;-A�~ �i���x��e�eک�������3T^ı9<��,X��Y �L�>Dw��߫~���[�T�����4��,e1�h}Y�F<��E��GTڋ�����2��LBX?N��ɴW����V
�FJ�EJ%�Q��Rh&���v�v�`'�d������;���	G�"�7ˆq��yY�𻍰��4�X�/0�-`b��Ö+��As^��faR�2��=7 ����WC_B�d"6-R�1��ڗd�9��sb����o��W�Q�Rj{Q9�ɭe��t�_T�4��Z�'U�o�P�*L��d�H����������i_h��Jio��(��#9ȔR������-8���J��j��J$Rv �Y�|F���u�0ZΪɿ�%(�j����9�g��Bn�${T��C�R�3�]��|Ѧ�ֻbI8��u��w�Up9��V2i�U����b�wQ Ko�H��+�n���ZN#�|
��W��km�2�{�"����L5�SZ�tF
�[z��T6>�;}�Ά�Y�xwa�XƸ��]�V����%����u;K�<9`�z�O>g�S΢��{yk��'��_�� lۺ���ٺS�W�E�Im�6��'��:�9�`���L�v�����Kҷ��,�ʓ�I������H��[@���}��}U��{���Ƚ��ʯ�_�۾����P�#���XK���\�Ȟ���Z�)IQSJ�V��5ܧ��?��B���6���t%��q�G�R�Q��@���HZ���
l��F�p�_�+.ͧ�����KE?߱�	� 1��Zg����}!1��t'�{Ԁ��׽�A֗]g[S˯Q�b�O(T��5���g��F���6��_��0�3O{��H�l�=���x����E�hB�-��}�Bub]�4�^��^�SZ�	_Cp���~��kw���i���[U`���K�\�,Vy�����!����j���E��*�T8���Qw�BY����x����s4p�m�_QD�1�ք=��/Ҕ-�Z��x9�O�H��|���ԙc�����Sp
���mu��(�`6f=���z"[��l�=�έc�;�:ֽw�/,�ֈ��T�h;c��>E�e�4E�1��O�1��3b1,Z�$U���:j
�j7�*���xL
{��sV+�!�tU2�w�m��&3E�q�̅�~54��:����V����d���$���,X�Z;����b]3:EH?7��a�yM�q��$�&d��ی���mVz8Xt(wL�0o'_��� td)��]�z��HM6V&�>�m�K��O�����T��ޮ���������ݺ	B�8��9*�#��Y�
����?;��I(�Z��u����\�,����f�kuh���t������_��� ���EH�k�X{s��ੁa��s�ED���9��aJ���h�1��ѵ�N�-��wjb�=nV�XD$�߷u�2h�o-�&�Zs`Sڴ�5�σ����w�6&y��I�gVDc?����dƕ� =�*=��� �G�bl�w��1�M?�{��f�䩠�!MR?��O۞��Ue���SH�
�h���/vCC�X�=2|R�4̸�`l��C �U���̷�$0.ށj	 �6���Ѥ��?m��ޏ��GI���W��j�KS*;�gC&���sR��
��s�?�U"v1��,?Td�-�h	�>ވ�_�u6{�0J)K[CJ%d���5	5(��C���� �-�$k@�������Л4W&-�6,x�{h����t��)٠M?��F9��ۇaj�5�Ah�Mg��l���wÿnx�� L��݇����i/Zx�q���g`�V'U�����#N��~+��=P�hʷU�q����t��5'��V� ��$��+{yG��I��#����U��PBX�[Q}h�=����a���+�h��nh�!�/Cr�;�WH�.wX�jW*�.��U�"�g���R�ֲSV�����e�{Jr��t��*g�ɎޮfBZ��8���U����r���K6_70$�0��1�����B�,H��k�h ���\<[����O��B�
A�-
�4���3K\S�}*(�ll�6&~/�T�~-��9^���[V}H��e]@���(�$]}������k=<t���(m�~Wu����6�b�����ͮll�)R6�zM��>�۔=tg�͈R�W��k�X,.��h���ƕ&3��|rl.w���������V���?��2����X��.�wu?lӡ�9}J���Ng!���g|R�����B:����a\����9�Q� ��5�O��d�@	a�5������FJ�f~���Q�n� ��Hg)����ЩWP�I17`K�h�a�&��0������N� �͆}�5J.��N0 b;+��_YͶ���z�5 jN���rX[���zH~U����x�BYw,��R�?g��\�>��D\�Jd��w�"�|1���D+<�	����L�̪ҳ��P�I� �gY���o�+hX�+�Rp��g�d� �v�(�H6�e!Y�6g��-�V���m��y�}	�QQ"�����M^?��' �*����~��ѓ�F��e�!�y,�����kf�⶷�%�z�jc G�E�s�q�M_����g���8	-ďyu����9��j���C��a�����bgy*���5�fs�s,�u3�,����~)Ųս�Z�i	��$��h�|��#"dhz4���_�N~\3�p�
��|�ʴ�讒W��&�d�l��L��[�9��Li[�,$2����26��U��B� m����x�@�ޞ�%|�8��3?��*���r�x��P��X�4�� P�Zv�W��*�/��A~��[�4���J�g>���c�,��e.(y*2f,n��΄BQ �ϴ��#K�%��t��6t$%���O�V�@W��$#�}��*�E3�-���tUR�rC�D���۔F��N��
I�3�K^��KV�s��(d�o���b�ʢr��Z�Ou�wwʣg�q��<c��ڡW���:�d�ch����xuHW��mL_�_"��o�:T;�9`���&-p�*����(�,����*[����^Ւ;-��=l�>��l�F��HY�P�bi��/i(���őiޯ*@%3[q&e�A��T������r�㓹�,���+�]�GR(6���M�\��~�y��_v;�'�F`5\��G�WGE�v�H(%� -�!)��%�ݍ���twIHw��0t7��y����}����k�w�g�yώg?�����X!�Py�S7��&�iCm�6OJ ���P����Mr��J�7T�`rN_l�.��w��7��w4�NT�lϫ�t��5�w΅��SF��KF��<���xkNF��%�q���N��'�N��R�.�jX�p��6�2����+YT���ޢm�Ҧ�In�w��\��3�Z�&Ư
��1��^1X���d\RJ��V���̻PB�U7Ѡ��x5��8�q{�@�X=.P�C����~)���zI8x"�+m6f3��p��8��o�2�'J%���6��ҕk�HnTshOa]j��&$ޔ�)�΋�E$7�{5�LGGӧ���7k��VK( �s�~�����Jt���Xu��<��A�7����9�� �㒐w�����"N8%&�C��#΢�	��x�YIx�!�F���;{[�*�ƀG�_�Jbs��1�J_1��s�ا��\�xm��Y�=n>��M��$7�w��J~|ǥ0W��B�8�D��rP4;	��ꝟ���G냳���w�&=���<"��*�sb(��!�6�O'�F�4tiX�e�ĞqWƴw�ޫ_����Xn?e�2�\�����8��[Zz�'N �H(��k��D��� ۓ,{U���7����]oH��J{eU~��.I��r��,v�fF�awt
 ^d��8�~�*��y�d�o�b�D�v��������2R@�7�ʘz�]h�#=���Qk�{�x��sk��`&.�{�љ|��[�vt:�}�d*b}���'0�}sAvջ�c�Քк�J7 ��M�&�k�d� 7��|�~�	��i�I`��<�+�敮��hI�kު@#��a�d�hs#;.j����Ķ�֍H�Mm��ͧ��Zѧ�pX+��=f�t��T�?��U�)������!8M	���5��d�5�Y]mK3���:��/�i-e����j5�6�6}W?��H�^���p��#U�B����x��[3T���1�z7=�/E�_�ބ�}�柳4�ggb��r(��*�[g@BUHP�h)��dp�TE�0�$|k��5��^����YD�YęZ)�îi]�B�@0��d��t��Pwvkw�T���$σ#:����c�@* �S���D���2�If)�W,Z�m�iU�~!��{�� ��~��}Ů#G�/Y�2�J�L�SE�U1zݵl?޲i��eD��m��J�W�e{Dz}>��ATb����HU��@,�q��L�FTH�S���`�O?]��Pt��7s��⇉.����x[�7m��]��@w���3d�A��7s����`/	�w��z��5�\ԞF�9�g�ͽ��:_�5P��Hפ��J���ر�a��e3� P��3���5��cS�_�p\ժ����#��Ml�\�6�m�
&�K��J])6ՀY��괙��$L��R{���z5?�=�R��*������o�vKC�]nB�RzK3��"U�Ь�+��L̖����ɻ�nm�w�IK�̄w]��ˤ�4qƒ\��@��x�_)�h��	�YF�\��d¦&h*�\�r_L<5{�h�|��U��r��ΪNC�n#��v'���j��v���c(i�69i�U�J���MmE��]�g��H:���2�`Q1)K+{(�,��p�KH�>	�]H ~8�w#q�f��_�6��ܒ����Z�	N�c�W��@K�nV�E�=�һ1Y�d;#s�d,Eqxn�i���4������i�
Qˈ*V)�#�]�7+�l�D��������Ǫ'&�_'grj�%�����s�T���uX�[X�u1���:j��TK��5)��7$r*&�{���q���q�!�G5����E����gK�,U�����2񉄿�#zf
�*��3�;`�fQ E��p.�y}�o:���%?���yd�W�ަ�l���ꥈ$:��V�MU�����s�v`w>'駝e��y�.<�f��#c*������/m�8����v骴��	��v����6+'�� |(�&������?}39�l�mǫx�������Ԃ�������q��_��	=�)^�|�~�v���D�J����>WDL���\�����wg�+�U��a�}s�Ic�;�8S%�Uar6���f���[O^��y�e�9b���[I�/�[=�}����9Dɤ1�,I������Pe@�����p���+���/Ihq�	~W��`���������7]6ϱ�WMZr�'�.���w*���W�Z�[�pO(50��ؙ��v���эz1�
 ��*���{'�@���<~z~=�b]`7~Y
P!*����T�)0ET��њ^�Dr��D,�+��>��5���g3t;b>�$:������{/\_:�
�z�"�����s�E[�E�G��q����e��ާ�(;�ƥ��k��72�=�4.��L���+��<����9e�[�k	020�'�2��F#G�A.Ǧ�/�.
�M��R��ʛ�Iz"x����k� nB`R��\��g��K>l��j�c��04-�����5V*����
d	r7�Ā}�u߂����ٝi��VXo#����l���;�X-j	�i�?9����
9}A�����͌b^` �ھU?�x-m�@�p'7y8���|����C�k�q�!��{���]p��u��ǻ�l�V�e��v�x��j._g2���yl�2��+e�4����V��6+6r��Ȋ}.vY2�Y�|\�����t�$��\����q7w	�Ш����W�
J��nBdKC{��E�e����1��E���$�i���I�F�|��+���e�N�7�#x�|�,N;���.��W���9�����C����U� ��	�˨�f��
�R����!u����������2�*e��k���]�bV)�䦞:=�P��ݛ-�?ζt;o����wX4���to�Ǉ���mg�7���ט3i�7
CA1!<�����*�^P2ڗ�UY��H�[A��i>[r`���O�
i{3²=˫z&oO�SI��X���]B���ɡI�X
�J�E��R�_�E���F5�J�~F^U"��`���Иo�FUS0��R�TZ]�r��+�%_Z�{�% �4�*d���B4�X�;��N��w%���U"n��-���Ƃ��Q5"�*7Y����FvϿ"Lʸ�$z~�
�M3ߩgj�t��9=J�zO���s<ws��y��Gô�>��L�Z�FY�������]��w�A����2WM(���(&Sê�E�PP�#{~��k�����u�b/��旲�y��ԏ���}u-��sg�*-�	��>2Y�u�6��
�l ��Ij?w��r��g��{�J�=g���X�n/y�&O�B�xW����R�WLYe�&s̑ޫY�;K�0�w�*f��E������ܷ?�%j[�ϙ�[��na}�Q~�[���wӆl�zb��"z�Xu�h����2���.J:��,aX�0PPF|<{�W�����Lin���Z�Nݟ{�cl���g'�	���������k4'\��c�E�%���T���:ܾbUق�
�OKk�m�Kk������W�?�I���7A���%c�<x��&����:�n�X�{���>��px�OK�Vw��w�c#��F���ꃗ���_�o��w�	N�wN�ⷁ_�����}��Sk��5�ӌL㷎Е�4X�R*ӆU��8�1��A7��*[_(�n�������ɪ�P˩-7��f�ܸN��9�7��Յ�{,L	zؿ�e�~b�{}5&�����ҕ����0}!S��*�^�=�ǟ�ء�L��<m��Ti���^���~*�Q6/^�\�|x~ۚ�0�xe�^U�f{i7]�KKp�I���[L \}�3u�"�<�~����>$�؎}�E�h�}�\�5��Qf��q4W��O��/��j����L���ớ���W,W3@ჴ�jޝ�y�|U�uF�:L�I�س�m�;����d���!{[{Z ���0��a�Yj���X�e�\�d`�u�7�R��c(��p$���w'V����Z����l�h7-��jlh5P=.R�	,���Sv͗�K&2�A�g{-�n��BE`��\hµ����c�����ө?6[��|7�i�m��4<y?b��w�r�G�	�k	BA9֦�7�F%5���i>w2@W�6n����۾p&�o�X�>�e�fla�"0w���zc��!�ԫν��e	ۨ1�r���VQKG /�����#��4��P��i[U��Z�( ��|� �u��J��a��F�A�9��2����}sW��^ D�ppTƇ'�g�לf����x�"=˙�Ј�}8�8nK���<w�(E��<:�G�G��rH��/�9\�q�e=�qp�`|z	Z7 ���d���4�<�@��ڲx2�[|�|�!��No�X/~�S��N奥�s��F���a���Y����˜9'~(�aW�:��M ܩ%�x�a�ʹ�Ԝ��h�PQB��Y:�5i���;��M�ow�z��'������܌���b+�K�z�µ#hc ;ܐ���t�>��t�V��g�W��^ڀ	��`q��3N��a��g��f�~/�$�u��%�T0V�zo_W7Q΂A�v�{�����2�廲W��w~�D�H�e�O���B��{(W(��,�~��u�@\q��]�^�qi�|�Υ�"�nBf���@z�|�W����! ـ;F�DM����ID�k�;Q$6Z7+� 4�u�8\O |����ۿwX��?k�A������O0�����=�ొC�{81L����;Cל�Z=��e��( 2��k��e�_�5�����v�v��,�WH+�]B78��|"��3'�9�c�ْ��)Y��. �|�'.�����cu09�U�C��<�A�Y�����VO��?��jzt
����R@sK��F��r>��K�R�6b@��๡���C" c�̅��!���2�y`'S3S�]�y�c<�L!�>�+O�����l��,fA/����?��I��η�=����jұg�r�r�'�z�ȳQ=��V�G�Л 2?���/,v_�����}UC�y�HmcO2D�Ѩ�k�v3@
��O4��� �}��PI�I��}	FPC&�P!�޲��؋��_���y�_zʨ$pT[���Js'���J�xi(H�2`�b���b���e�����K5g�@�z�հ[�ǒ�۽���3鈭N�v���>�UQm���@����ȑW��M����Zo��0��Y!2��O�Ս�y	Hj�+�C7�ط����y���nZ�D�����Pp� ����(j0���zߓGt�AI�Qv�Ƨf�Y O/���ʯ��m~�?�S��'��A���<�)����_�����G4�[ô�6>L�f�,���ޡĲ��n��B��$,毄m�����y��[f���13��0��Y:�)��P��I�BTA˦3���m�����Ό'\C�aZb�7'�9��6���^C�a�z�<�B��A�Fb�B�+]k�"�#D| *��������z�4g�E �XG68;����+Hf��\-����!�0���roW����%g꨽ ���[��}]�3�/郶}-!���Ű78��|������lQ�N��E����9�y'�e;d,��0����r68ȸ�}��l�I��l�A�������V��b���8�;o���E��b	O��SQ!Oٰ�v���B�(�������J5�@%E"fq�R�6D
���3WkrQ���4ǋs����i���=��\4���6+'�}��~*�l���l�}:��<��TlR�as�CyC�1u2@�_+���Y���p;_a�d{G�%��ws�I���B�;t^�/���y�D�+3�J|�����ݞ��P����k����xX��!de���~�rx�������xF9�����m5�i�q�e(?0�N��w��5�B�F�VO�_rj��s�zRH�nl�)m��N�m�]��л ��\G]lJ��3�-!�G��]!��E����O���ע�$�l��"u}��ȟ��K���ݗC������VK�^S&���u�z'�C|���TF8�xn��*��@"�#��si'�_��EIQ��rM��MqX�M�.xec%D����=���	��#�@��!�f	�1LB��&���������D6W6P�[�%n �@�AR����R�'9%�W<(}��X�.f�Վ@4V�p���i�n�cI��k�:�A4��/�{,>�F���SH�����:R��S�W����pB�D�s���>5���[DH��{!W���p�h[s�_ �H3#%x@r~�H�H�`qRV�����D�\(��i�<�I�揇#��8�yH�"�{A�R�ey��ݳ���*������G��{
/���ڶ��y��D-�*�?P�������Y�D{[c(^�hhRY��;3�]�%�1�=�,�z�Gym�摤&ȿ���>���kǂa2�o�������_?�[3(��?*�5܀*��o��䭙�/s�f�l����0����$t�$	���'q7yiF��l���<��^n_�&P=`�;�ӟ�(b��W�h7�)z�����95�� װ�xxw��7~�i�1���D�'�T�EO|D��qy�`6�>�.������P���q��f$�bt����#��\RDg�T�0	�����í��}x�	���&��d�'�޴��c�H<{���e���M�4�j�մ��*N���s����u���.�+��mT�S,��Cc^ɖIJ�j&�I��⧘i�K�g��Y��F�N�}s��Q:�W�ELo#�F����$�y��	,�<����������q#5���PZ��W����C��iY6Yn��7X�/<�"���CD,մ9�H��)����Ip�	�����0,In�_��������ߠ�'}��E�*��8D�����L�/�G�����1�_F��ݡ!����6��SB�_7����?�}}����c���J�|7Qd?��T2�g�E���z���Jd�ma�TA��JzE�럨'��͹?��-K�T����o��L��� � f�p��ۊ�|�\�y�<�
4�k{�@������7_����RN�_�{�,n�ED��6:�$y�����Ab�Fr��L�/��I��V>�:	B���Sj��)��2(�#v~&W6O��nE�g�^��ҡ��3��l��^|V���?q�%eR�����f$����M"�qЃ<a���(�G?���5�p�֛�}��lL��Jk�C܁6��~OA��h�!����q���yI�LsE���e��G���ڂE��@D2�����&u��C�]����M���iҸ�:L��r�>�ѐo�JL���.-�����D�a>���̊�3���ZO�X��鵡�r�oʞ�K�������J�H�g�*y�~)�|��"b"��g&��v��ݸ�Wg�R�A�h�'ʪ>��cE���P���^���9�S}�I0�k����!pn�R�B`m���#��3/�྽��[�z^���Ǆ� uQ����p��lvkDuR~�F�!�ʃb�ҟ�g��G��q�νr9|1<�t����.qc><��AL0�����ŗ��+��:�w:�r	�c��~�\�/���5��	������)��U�^ө��({�#���6�J���apsh��=��'��r�r��s�MA���K���L%��w����PH�^�H�ܝ��=)ې�J��[lD���];r$����rg�cft��K��ފ���?���;��$|����Ҥ��>��H/�QS�P�U����fkD1���s/M�#����T �%�����^��A{[�E�#�IH
�!l�K��#���Kt��B�����Ʉ��,_��|o������l��"c�Ly9��	�ɰ�����nk{I�9}��M�����&���ߴ�iW_�~|=��B{/,DV����&g�7paw5j�sUy��#�Rn�p�[+�o�e����ٛdCu\��L�4��D���nc����D�U��,XQ� �p�R���5��Ɉ��>d�a%Δz�]���c[/ޣ��E����g�n��q2��%��eg�ޛ�ʛŴn?z� �o۷��~�s�dU�`fRF��<3�r���g������X�=�c)��Ta��W�����L�i:ޅE��z{p-��^��nZ78�o.��ak󬯕�N�{�]QG�5;�pf�T�ʅ�?��}6���~��#��U`$mˬ�G�;B>�<:� i�<��i�0k�w���6�%�h�w6HܪT��)�
�A`�7�$z8�%1���� '�������D�����Q����Y_\㺕kw��6��BQ�y�O����bv�6�ϣ��H�㇟vg�-�x"�\�\��h�1j枘�D\N�M�6ZД�rV^��s���V�zF��ݚ�"���(ʺЏ����ȸv����C������ 꽻�,�wu>���Q$i�:�>��Q�������yU4�OY��	~�Z;�� Ä�iN���e~��� J�(X��1�E���+��nI�T�����i��cv�O����'QYG���ڍ���r	��u¶c,��g�a<It����i�W��%i6V�%��!�H�iÉ�q�/��͉8�"�fs�&H(I׺t��H���E�b��h���8�X[�KD"^�o�$IC����7O�X��c�\��y�ˬ�XCiJ0��Ɉm�O�j���X�Μ�����n���$)�!�F-�}���$�Ǌ���taa��������k��ٺ�^\�k�c�uհ|_;�2݆=�(�nY+ߵw,�����Q�ѩ3�6��=Rѣ	�P�
�fDT���z�L�w�R+��K�3���ˉ��6��I���y��\���,:��*�Sw�E$�t���dE6m{�K�Kwp��2�3�������x��a��rx�E�K���g���*���C.!%����#�����؃���,�G,8{!�.���ؒ*�{О�\�6�q!K?Yn����Qg{�d;�̹ޓ1�W�݆��g�٤z֮�h�q�3���4x^�}�]�x�]�Z�\u����®�r��u| ~���m}��u!:������po�&$��A�0�"�HKvi���![6kMS�WL
��楳����;�����͡%�_Lw�O�/7U0p%��t_��+��g&�%��V�М���o
�v�jMϏt�� �۟�\h��g�ܟ��E���������ڔ%콵.�߫�
+4�0��B��tD� .H �C�-�/j�TT������	����m�(֐U��R��8��D���g��c^�9T�n*֕�Z�aćS`D%0��q�;=�Kn����	�` (ܮ^��靴}�OȺC��\��L���8I�����!5���Q������Z�eS�-�dmUT��l#"R���iO��g�l.Ǜ�FS*�nh��̈8���N���fH�$�k����u�j��K���y��Yx�<���uw̠G�ڴZ�C%9��5�Zf����g��Z��s����^��+���R�wb~�6X�]���F��<񃁣g�������Y�d���_}|H����$Y
fZ�.����$�� ��Ҝ�Ѥ)�D>�F�ﰬ燊�kOc!���m�k/:e#3�:�4�m/��#o��65��DΚW��:�;M�w�է'W%MuV��_���=KYcW��5��*� �Gv�@c�sprn���(�u�  o0|�[Λ�7c��AF��Dv��0�2����1�#�w���[�҃^�C�U!�3�\���u�
��>�~ λ�_�z,�ɧ��F�'����v�����L��8�	_�~q��T��/[j��4S^<�������(�;e0�MM��ޕ�P��1%šM�T�E[�fC8P��J�2�Z�c�jP������"Iz7X���.�zMT^E��\M()�o���S����E�����ӷu�N=$�ޚ���#E���!�������4#z��⃌��_��p���%��z�Y.�D�(V�H�g.�}��cw]���p�I���4��D�ř6s�����6�[�O�4�<y�eW���^�.R6��^�����e�
��` �t'����';-�且񵼇N�zB@%QŲ8���tM�2���0�����W����Z�KhF��|����O�`��j�5�J�q�X��X������o/���Y9 �8=����u-���p��w�ą�Xhx)yo�YO���f�����&5ux��k؝[����#(;ۚ�:j�v(1��G��r}��we���g���e���D�/�vW�Xj���e"��f��c=�Nc���P_��n��~ =����(�v7����y"<���f%�_���D���4�q)u��Q��;����¬5g
f(����ӠԎ֩9��Խo��¼I$��g�A�8��+M��0�!���ˎ���-�C�@5���F޻�5-"s��°�xjZ��c���DW�DU��H�o�V�����C�K�ݞ��*�Y7�H�GF�S,	ӻa ���/��x����J�S <"�|��O	Bw��us�)0�i�8i�������ϛ�~/U�w^�nY��>"f���/�_���5+S��KHh�;�Nv\4�c���i}e�Le0���M�"Bod��Of���N��H���9���z��hAH4Zlf�RY?�N��>M �������J���~#Q8����l1C�O��t)|�>~׆�T�GWy�UUή��ʋ�-���T���ιϵ �[���� ᠞Z�+�abȚ
�ㄲt-X�hb�{��~DF��Ӆ�v���%u�	WQ/��`��W����!�$�kȺ�B���{��������=
�Ø%~0�; ��ՀZ��]�BB`{�b�I,�ݬ�ez�����>�R=��E��Q��Jy6�c� uZ���C�oe�����!�35M6}^(����}��F�ks�{��혦?SZ����_�0�~P�c;��H�y�ڧ��aJH�"��� Z����R�a��<B)}�����j�*1�)&Do��W$f+���.U���4�{F� ��l\vL{4�����l�3�+�PӁ���*l��Eܐ�$�n"�7kmpY�+��Ys�^8�j�f�w��ǡq�����X��s@W4����`���		2��5k'��ڢ�"le��w/�a��V�S�8*�c��^G�ݤq�h��R�1��΄b���#�{U�B�b+[�����y�x�\oR�td����,�I�a���w�>����t��Ƽ=��Y?N������������[ż�s��ʺJ����h���.q[���M2`�Bi#�W�ג]l���:�y+��wU?��Z�H�~t���^o�g��S��I�L�<�DHV������%;�5�/koz��`"�.i{����@��Rc�9u���@��\7E�~YE��*,I_s���$w�.-�r���W7���5�۩S�M����*eLg����h�h���b����b`�,���;ݎ�D(]��(9�|�� �O|��H�݂��O�#�~�[mG?��5�NZxۻ*[(ޣI�ȱ`@����G�^�t+�Ȣ9?��Z��PJd1�)MR�Iv�.7 /G��Q�Y�1}'*�VXu���夞k����/��	1FL\�l��kFҧ����_#����M� ��Ѿ�_V"=��9F%�����sT�W�cz�7Ak@0�E�� !���xqփ����F�d~ˑ\�^�!P�X����q'
(���o��S#�#"W��n�ZF���+ԥ&x��z�\xԁ�hF��.��e��2+�N����m��g��qEW�2�2.j���!v��c<�aWbw�(�HX��I�i<"�:I���&�7������U���]�QIVQ��N���'���"�.���kv��Y�J؇�bF�֧��h��T��ϱ",�h�� U����Q+�M�,j�߾�:��80��Pf�W�}����؃z�.����S�26׍_�J�X��۷VK8��x�����;�ah+������z���]��A�g�ڽQ�x�
]����|��u[0wz�SQ9p�w�7���T��O�8������C/+�:\Σءu�Ϡ&�s���yxd�6([Q�oZ���ĺk�d�d�e��G�	��6߫]!c:1��6����Q>5��+��5�u-�D�"�r�r	4����EAW4�u�I�_�/�]ׁ���L��l96mq����bc��u,�t.{i�*ֶ�`hT$"�D[�o皦9����绢c�T\`I�N��asm�Z �����{\�����'��DS�bԵ�9��5��\w\�C>yp��b�Cf����W@̪���P�^9ΐ�!1r�e�!� �4EŃ@�NZل~�����|����x=wDַ�'kC���e�b�Ϯ=!��q�Ux3����5HYF���Q�A�mfH^�
�M���P ��7�,fk�1��>�N�J�����&�	a!11
R)1��Y���º����N���>���`��5n��-X����������hXgG.J|�s.,T��8Z������ۿy���B]���o�ȈsZ�V1������}��A|?��BY��U�4�40��`c�&ӂ7:Ѥ�"�'k\Mff���#�����Ӥ�v��*1�:゜B��������F���4*(��~��F���$0 BJ���[���.�)�9S�ތJZ!�A��"@��}�����noپ._�Y���H<"_�ҳޚ�X���"�9S����I����:�ʲ�A�X9����a�c�7[3Snl�jW�����4�W�"�"��k�I��Ϯ��8�N��9n��oq�.�3��3MBa̟���ѦKF,�=�aZ�r52��fR`�d0EY������6HN�ڱ��,�V�!�rr�헒XUs��'-y��8۪aRto��zk��+�g�H���?ߐ v��	~��@��A��<C^�4��ĄpQ�S��R�E�v@�<��B��>�U�ry�������WMO��3�K�я
 �߆�nV���"���7�ǳ<7�d����nA� 9���p��@��bTo�<d�IP�*F�[t������hL����-X��R���؉5j��3O ���~�����o�%58F���
M�2��X���:�|�`�u�	��ۺg�s�ٖ�%)��t;ihZ\.�Pݮ0QTW�YS���/4��)��J��F�{��8G�c�G͡�d��,A���\W̉�z���˟l>�fɵN�V(+�V��E����٦K`-�!�pG��OFSK,��?���l�l�y����dK����0��!��Vܘ��5�ymC7��Fs�r�>̓�w�AXq|�S^UiÑ��=�|�{��Ɠ���R����	k����S���|Ѓ�J-+�xޕ��.��*��0�k�Fz���S�B+q�#��.c�?w��q�Z'��C�}<N����V%���q"��Rio����mI[tˉтej,�&&�w�T,���L��O5�H�3���X��,�qT�B�@&0���t��9�����ڼ͈i
{nT��-���GWBS�gWt-���-v=�t��x�t�S�C�D׬�^��ܽmۿ����}��zt���Lg��۷u��6��x/���ì��IҞl;�֘!NU;~��/��*%��7FE�t#�~���!�/�6_�ڭ��5F�&>��'����ir<C��>�]!�0��I��O�b2L�Y���������k���z�����.E����5|AŮ��U/E�T�a_rU��e}h��Za��Pf�M��q�L����RI^���s!Z��<����_2_���'���#s� ) �-�`�nP�7%/yc9�	�U��㽧�7��F(��Z�	0f�~=5�����JY9@�]� S|�~�i����1`����|*�%��J�`g���d1��r<�+=C�	��N�s�SM?0�;$�[7w��ƕ����56^B�
~c�F��4�ҷ��aCh�r���iꥌ3���;q��"K��b�>"�XE����@G�GB܌�?�4�@�T[���W�W{�K5��-����$�����&�q�X|b>W3����x��Q~
Z�Z�n���~eO�fJ��b��;��|.=6�n��=���^�*�m��睌�� �J0#�Jyt�B��˚X_ټq��]>���n�q�u�vq�p��j��M�޷~�˩�~AB��$À���L�^h���]($,��3�>�tF��t�����d-�>�����(���ϛF���е�i.w���8��	��Kl̑�)��?N��7�جt�L1H�T�0���_��N�I���}˜��ꇯ�(,��Yq9ZN��5��%���?&cر}��E��.*,ܥ�h��+�P�ov��O��|�2QM�����o2��#��hU4�~Y�J<tI׋Yڟ�|���!�6�r	�NS{�먂e���c�K�b�|v�ۿ�J?�WS0���1*���!ո��`� ���.��ZM�2�6XںI�!��/OĶM6�P�`�l�#���9qa�5q�����Zz��L��;_�4G"y2o��.��'Ϟ�c`(��c��W��I�R���T#���ᰝ�s<�p��ާ�u��c<dp�#�u���u[��KR���B0���OW`b��/x�7|���kO���SH�+S�z_��M(��fd����]�i9�9ps@���rA���E����-���a��y��U�F��ޯ.$Mӂ�c��Uc�O+�"0���(���K�s�[H��; �"m��띵Ɯq��A7i�y�g<�ؾ~�c�I�����{�v���D~YZ��D�g'�+Á��KmCG0E��E~¡O�?Pax�l�[�>Mt�sU��?<�E�j�u���x�61�����8�ԫ_�6Ӊ]�����w��:(*)OBi�(�F�m�B��;LoE��c�q�g	�)Y	p�R2ߖ�W�Z�X
���k)Ss�z�uG�K��燌�O�����((�q�@$�������t�g��`��5�Ǩ�h�Kl��M��N�'��a�{���+��1����=�&|X_�]�7u�~'v6Z}OU	�U>wh"����Ӧ�.�C~��Fɍ4]P�7A�Ute:qY��\2(ڠu�����"H;?.��Gr�U���|�֚�?�}�nz�� �� ӛ};>���pe�'�s^K6jh�9�rN��S�WW��Á�O?̘������5�Bx����<>|����k���ҡw����&�q�����?�?X�rb~���&cc��-aP�n4�p��XN�.�t�Q��)|�N@�����Zo0���#�:��#�y����\a3������,�<<ǎNr�A1_	N\g'K���o?�X_�	�'bkI�|�U!'���P���(��$����@pƕO��44�m�ESn:��r+��{����L903�HjEG���)�W��].7��/�>������K}5,�t��Ų�V⍗@[K�坩V�����������T��\�����>�c��`�R�v�ŃK�@�d�8L^�v>�OS�/PQgd�cV��ރ�#�/Mx��=���$3H�.���Q�Q��&�<�"]]6?�����������I#E%�Us�E ���`�KW���um�]��S�o�`C�&7W���קx�&@�"u�q)�ה���c=���˖C�]��S����IWc�_Πl�@�V����V��1��vg�w$ �r����np:	����Ƚ|��/4��[���9���7p�\���~�t5� �]]�iZC��}� ո`�"7f��PY��>X�<���,�!%�;��H� ؖ���m����Oz�N��:rK|wP�,��X�5N¬��Os�B���MM)A�W�Y��ED�"��gE�=9��پj��p����R���'�����q�B�:���߷���DW�ob�ۤ���g�˖��=?�j�6E��ļ���g�!��z�C�i*#Ď��I�x��qN�1��@�������ʌ���s���؂�I�I�<k?��Ul!�(���	�O;��c��$^%j�}���M0g4��f�w{��T� ����+τ@�![�E�I�sJyl|K���Ҝ���Ȇ�~)%(�j%Z���������~Yh,q��`L��E.v�����vRGK�xc�P������
i7ב&vU�u��o�Z7솒F�1@7�}�.����f4D�W,4�:�1��y��u�K�9���x��~���&xG�@3,��u�g*.����M,����j�m���j|Y���/���� ^�_v�
{�	^&.@g��h WQ���p���|�y����MD��++�a`���ѹ.?:h�0���Cu�?t�@�}��`k�'A��v�6���XLoėޜ Z �G�4/�rA��!Z�m��j1M������_ߖ�_?ɱsmUCK�#i�lX%�|' 3C/QtRI�=�Q�#ȫ�c���-1�&���}��#2���Lɴ�����P����z靰AN��\���/��|2�G=���۾h]�bz� w!t��'9���i��㝲��v#N�����2���xNv̐E\�K��uk���z��Feث;����oPr��7�8���!^N��>@�����H��V*�
xᕬq�l2l�$I�ñC�%��+��ܭ_Џed1I��%��=w�+��8b�F2QS뭫�NN�'t�K�;oJ��e!'�ڽ��$�݌e�A�R���Ʈ%�<��{FC2��{*�"����dM�_�����k-q�0k(���Q��)b������Ɏ�G�`},5�@���JV����ᎀ�:�4ֆ��a�G��[��xsC.��:��$����,�:��5�3Hf�d�LS��DJ���x�+!��޼��!&f�][K���P��ܜ)hck�!V�n��}U<�B/,��n�xF�p|%>}����H;�-�˦>ۨ�Ւ��z�;ĲQuaVF�}J��>i���;�	�2rP�?d}T�o�� �Ej  %]��K�[��ctJ#$�K@)��I�]������?��s8�1���}�s���w������˽Mre*}����d�|��r����{��I�+%-��kS��*4Q�ԇw�8����K0�f��܄'��_g���y6|�03���֜E>�иf��!���"
�Dɇ��6��6d���������E�˔��_��T���ıh�0C�e{<┡f)�8c'�*J	v
Ƅ�gY
K��9�偰_ܘ�xg/_/W+Y�=V�cj���G�f��n�ZS�'���IrP�=�an��/j�Hᵑ5����4�9�L�6����՞���<<����%c�=�)��K*��_��,�o��V�{!�y���şz(���4��*�|��
�����<�r�F�Ԭ_�d	����Z+�j|��}��/4=X QU#]�����+���4nL���8T�N_m�K�\ɰ4z���k��6U/��;�FeԊ�y��mH��E>F�|�5iO�3���m��z�{W���7!���Z����?	}%/���lQ�@1	ŭ/�kA��2P�S3�����hK�:zK8`�j��i�X�Iqy/�c�.�M��N����TR��%	v�N���k���H��/�|}�"�%Y��e��hY�,4��T���"Ù2�@9�M_nϡ���$@�F�Svk��81�h�28Ð���̨��}��Ċ��r��R��I;
�� ��m=QdO�:z��?��鮅=�m���%��-0�����ɏ�/¾����r]>yd �j���IL�%rr�?����ۃ`�t��\�Hl+�9����JkS�͟Кt��##H�jcs��<�h� [��3�5G�N{T���Hf�#y8u�*#��Z���w�H���xa��h�a>� ��q�~��E4��;}�Y�M`��_i���3#�Z?���ii3���=��e=��f�T'D�8ܰ���-Mt��g&i���]�����%'�w�``����������S��/z��<f���|u�}NG=��o*��Ë�5hX�jXz��ۿ:�o��M��E趞�����qH\�f�a�AG����칈�h5��}֐H|����Z]-'u�����T1�@Q�2]?�U��SxY��SY��_�����������������)~�l%�h�����\�\8� �͔t�f1����nj+(̔��ej�3����L�Ҁ��c�Z�8U{��}�t������L"�� s����׻ͷ� �+Vy?��2˶��$S|n%�]r7��-��ܒX,/:8��8�H�������\���l��:~<t7#�jPʂ $�_7s�3���u�����X��9���2��H�]pֵ%o��w(8�z.��x�GTtXIT��=�NucV�
C0��ߤ���(0�>l���SN��@���c>	U��g���?P���r�/���r�J��\ʃ���ձ�6�(N�B+<W���SSh�l�V�_ܿѿ�w���[M9cl��-�/^���MH
%�����Z����\�~����9N�3e��P�M
� _�v�z�k���J`��<�pC�;[k
ZGʞ�qo+��NEt�ї󀪩�r�vr�ɿ'bgϱ?��e$���ׅv����dlHx1E�f���n��ڹ�b�C��c�2 }m��986�����<��o�`����ezB��.]S�5��_�����L��EL#'ռ������}45vp��_9��w:�`����-�͏��P{�(�R�'Y���� +ۗ���j+Я"D�{�V��a�E�aԱQ�_���z|�u��7��V(N�ɞ���_>ό�R5aB��d<�a�\4�e0K�Ȍ�Ve+��W_�3dٿS�}��{�j�ςV��-j�$|��a��h��Qú?�˸��%E��H�R<p�f�!bRCSKZ��	):����m�-�kw�ՙ�n�˧*]�P�_���Ȟ���O�G�h�Y=:����~�ܯ�<o��-��NoA?�$�_Η���be����D-�Q�
�y�l�T��z�N��fv��Q�^��wu�?�D�E�=�rP��u�<nϧ�$Q�Չ�d׽ߕ���R{�~��S��jĻ}G����{��Gv7��Z���l��3
^u�/�44;�̓=W7@	D@� �a�=f�.��{|ׅ�*����})�J>ʲ���V\ߖ�9e T�7|0����@S�9V����v��Y�>g��A��0��=L��1O0MH�k�!h�l�e��{Ҟf�X�m��RONxg����oE�u��H���|S��-��k��n��q4S�w@�y�m�B^�!:���	.&E�����[;����|���,�צv�}��%_�����Q� �Ɉ�4��H�zg����~/x�\َ�J�F���U��aQ6��4��u���0�7oh�O��+8VL��P]n]��z I_��
�x|cH�B}�U�]X\�.kq�����`(��)����`?ӹ�ۨ�l(U�p��l�މ��%+L՘
��� V�I����8�������?
��"Z��T�*#N��r����Ũ��؈Un1��ϝ���7a��Ig�~��c��υ�[�:������q^���d����@�Lc�1-wp��}�MYo<��:EN�t[�ע&\=��_g��ć~g8��V��������m�d�`۾<���ѩ6�Y�k���}3d����]5��Ұ��q5�I���ou��a��z�½��:�zE^��Q�wݿ;m�9d�{�����H�3`��c��z]�_~�t$O��`�*krL�!���̴���ď�p�b�P�7)I�i\�̬Q9�R/z��/�?_T�� ��Rq�/h�e���'va]��@1`0�U��	��EvyJ�\�m+��t� gњ2X�0�Aֱ� Q/��+<օ�y� F1+������O΋��E���$��,?g�a����oL��P�W�/K�N!t[�b3V}��;�A�T\���e��=��x�$�Hoħa����=	+�.n��Ȕ�wĒ�V�o�R�@����2�UJ����շ�f�[�b6j<�����ċ�����E~]ڍ,�"	�n'־{�^��O٘Ln�Nݞk4�OfH�ٯ��{���G�<��5?Y�k��Z�C6�Ź�Ѽ���H���������F�s�r�~���l�k!g];w>�b���(�T���i)9�K��N�V��z������~��]�y3��ؽ�#�|�'�����{#Ī!8��ŧ����ژ�_}�����sGʰ!�Rg
�d�5!�#��uaAz�q���#5��%h�n���D����/95}�	��&�c���2{=�k_��Y��l��3������T7�E�;Ք>%���=���w��.Z���7G1�
g#��~w�� u߁ ��E.�Ղ@�n?���>��`����í������.G^*Z�az'=���/�ګ�wǞr7�� Q1��9��sh���0��L�#�c���Q�f����������SH@�;2 \��5^�B����K�ӟ:��^�fH/��Y~�;������}����i����F*eƈ�i^��������+���� �U����c���[@�o����"�Y��&z)/�bI����x*'&��R�b{���v~s���q�K�z���c�_?���d�Il�C���upx��=�՜/G��
����Vp��ȿ��ݵ�G�|�2���l�z.�ǻIr�����98Uq=y8�dl�'w�Q��1�V\�!�j&|���x�\9
��፟yŵ�R #��w�2��|:����"��x�h�]m((�
̎UM7�W��.B��G��L�`*4@�ޮ�3g^t�Y5��1�^?�'9Xh�x�VQӞ:���}�ނ�]����<έy��o����C�)��+穸q.�dDd�8���Fz�PFlo~�;nd=�l�]�(/[J�^�3��"0�7g	O�xZf�n�D�;��|�Z��=���ί�6e[`<v�Bn�}߭�"9KW yⳇW��|�x���$�Xd�*�W�.w�<���Y}�ռ�g�>��gEXb�;�g}�sA77�rR%�K��Ȉ���Bg�SWg.8�VΗyL�]|~�>����Gw�I<�cI)ض_�1
�P%S�}�nz��n�x��%�Fԏ�Mcd��#�l��&����I�I.C���=/��w���&/\a�^����	��{��h3�^LظC�q<��.���у��ˆ�h���|z��`�ܱ̬Ce�b6��x���.?oV�a4 A�ωT�_r�L�����soɠ'Q�%��*��̽�֎��5t��~�4Qݐ��<^L=#C����ư������ƍ�O��i�"��E��c����~uO^�*��f/����˻��V�㓢.�+s����	�4��p�������@�T��e����dj�3j ���BZɞڤ��Ƌl�v�b��\�wX=�{���v�yn�n(�?{xzrbog)X�Z��~%_ݱ��iѶ,QV}4��r����$��������i�;.���	�I�������ˌ�Z|���:�`%�g���["C�dJ&)"��Vf����?d�vv֖�Ձl��^ܗ���^����Ee��j�B�����{J����(G,PQhhu�%\�테��C����%8�P�V)�W"hSiR:��P��e�q�:�������V���u��)��t�K�I��E}�\\<[Ԃ����q��c�PU�XL�O�)��+
!���v����K�8�=t��֣���_)��~��^��<�{|^f�&�]0p�x?\3������|6<n��gN�LI�ܝ@�#H��^�d��g�c���v-��K*W�����`�������� �NY�@��T��\O���)���UVű#�T@��(�vP��C�:@�Ix�����*����]}��s���<�9Iͼ�4%:�MkF������-t%�M�a���d���w
�)/�K)� �t��*(����y.��rK,b�x���~a�s3^�:FV#dVD[[�=�s�������`�����q%K����O���u���L��j�_�_��[߽!F�Ƃ
v���o+n��E�P��v��v�Og��}C�!�V�z]Ȁ(�w�u�&�ep(�3F�����s��˟�� ����׽�F#euWf�.�<�G`m�3�S���8���I5}�O�����@6��Ys�j4���N��3�ģ�)x��W�z����}����<���K���ZG��Aқ����Q,y��3�Je���Z�]��n�F�Yh��q�������J(�?���D��U�y�A��b�Ae(�?���7Uʮ�6~N�-^�ų���k>f4n�Z-��\������M�J�߰�D6�v��{#y�G{�L|s��u��ͨ{ȳ�$�f^*+e�]��:~.�r;Y��d��z֖m��.�G霈�< �|��e�]�W/��r.%� �8�j�Kӎʿ�AX��/v⣲�\!���T�0?�h��c���2�۪���z=���RR͟��za��A �j���`��5����s��������J!4���B.�u[s�� ��g�o�n�a<y����_wǶMWo3���b��ٔ��q/�I��V=�b�J@��\�R\�y���^i�a�b�8��^�����NL��V�O�=��YF;P�W�'�?g-·'���N�>������;9�/��~�u�	���kZAq�^�h#�,nq|ɟ tu�]v�%&��l 
:6Nr!���iv]��Z(R���2M
[��D[$*W6t�2�`���>{J��%����U������*��;�pv�U.k]8�ƺ�ͤ��bu��UKPJ[V�F!>�C9�<$�>F�Vd�T"�#;�hD����Ƿ=������r]|"o�|�?g������f�/�ظ�z�O����o���q̜�ɳf�W�S��Xض�heLW�� �bd�������B�����v~�k�*�?N�E�7�*3�Z�qcK�0�2}�y���^�L�����c�<�	y;��3��>}�P��t��wЃ�q�$��*rM��9uT��4�_�������m�~����:��uݨ�Pzu����~uz�b%�%�«;Į��9���𳤇2�W���~�#Ձ�(�u�	�G�rw2X_{���PPi��<��a5���=��$��s��A%���֕�JD)_�Ơ��~Z��>8���2֍I�;F��U�T�Y��?��3_�1�˼���4�$���ڲ���:E+$�.kZ���̿8��� �$��I^��0Qf����.X���c�����wM�K��?L2���T����Ղ[-���2$P��PE�.�ׂ�j����殉'v�u���9l�]>�����Y[Ǫl�o�'?�������%,L�,0���
>,�.eIj����Q���~u���i�vx�C��BDRl����b��j) ���E@�6dҐ�K;U��U !�+D6j��. ����4;k�ȱ�3����~'&c� T�����:�CD����}��B2*�F�M��%p�]��h͈k�tsa/�<TD� �3Z(�spc�lHܐ�W�R/p^�ONNkhh�~(C����L�,Ɣ�#������o��}���]Q�`(�o�h����s�Ov�D�v��D0'���c^�1��Z�M��.�۩ˑ^K�j�6��bu�]�U j83�d[���5�yݰ~'3���b%|�j�Պ�UFJ�����������M�3Z29�����7������V��?���6o�4ɑ�rE ^tf@��C���J�kY�2q�
ʎ�Ao��a�b�N����6�BK�أ��}'w�x��I�t�Z١HӅ���y�J�y�����<��3����p��<� :t������_�k�͑�l���� O�Ok�\�8|��5���!q���<+���(�q�׿�(,�xF���n�F�fy�ݟ�@��z��Ƕ��@��S&�e���]o�j|~q��ʮ���;z���`�O�ᮕN)�+�#�m�m�pUT���~)o��BK��^!���a��W�1�,-�R���K�G�t8S�A�ո,p}[Q�+#"�~���t`{,>����_�L�����������3�&�1��k��0Q�9�ŰR�T"��o���� ����ث���ҽ��@)�7�X��\��Y�\�-�q�[�6)]�sE߃֢�C��m�D�E�FѾ���rc,���彞������9,�~��ڻ"!���t~.�`�<z=w?��I�FVTTg�6)��z���p��"�a7g������8�<y³|�b�6��y

TeB��JQ�Sq�!_���.zG`7BG/�����pz�K��x�Akbp8.^�����EJh����<�s�'#G3�T��U�y�}oa�{K�4���l*�n?�J�p�������^uXx����1��ֹ��9]Jm�U^�"=>}�Tھx�>@�M�Q��3{�T�%���
U���|T�#���򣺙-*��5�.�O٤����ȆAzmL\�&�
��bF)�0&��'.���B笩���4P6La훿j�>�U��Z@=����U�n���9eĎ��䢓M૱���*�Z��X�k����K���7���ٍ�/>1f����!"P��_��oj3(�`���.��	^��i/7�-���G����/�W�}��(��aM��>-�D��2h�ƏV���ʧ�@��t6n4x;�+r�``[���u5xY��kx" ��s���vs�ųz.��.��s�s㇑'�]�U��@��&݉'0��ǉ:C������`Pw�PЌ����h/w�a�vr%2��w���4�u��		����F�QK�@&��&�1�Ʋ�˓1���x�eAq��]��PL�~�SJA"Kd>~]li$k�~�&M�DB��l:қ���N����MG���H誘��;oJ�ۄ���+��m�2U?>��T�RPA)M����[��'�/��vqY���nС��aK�:c��������N���σ��]Z2"���
G�C�#�b��aP`�8N+�ڌ��B&)���t�yN'O���	t9�hP
6�L �+���5�l�jXً6�>�hG+�NFp����P���"���&Nv����V^�6�Ǻ�8�6�)j���>��(u�J�qv+��ۖ������k�a�z92\M���<��3m���K۴���T�(��a�j�/7��X�{~%#$��Ƒ�L���R}�if$(��[���+��\,u���� �[�;�G�v�P�|��"�H�?u������(�h8���B%���>��ײ������g��#z�����D0y��^)	u����f��+�К�B!R��nK򢧙y
�6��}�-$@mW�>���@7��`�B�U L=���S���e��I�g����H`E�����p��.śh/����`WӥhgP�h	�(cII5(�G&��H�̚�E�v� X���=�J��#`���/��K`j~"��ᕅw�7�y2�sҨ��j:��5"&t�������,h��g�VT}%��Z6r��X(�x�+̧��#�^!�t��	f� �yݤ5erpx�1��\=K�}� �Ψ"j���{�{��K'�XD1����+b�B�����߷R��Om�h/%ld~��4e[9������|�����`a+,?}�,�j�+�,��⌝���Lۄ��`��θ��z���S��ƶ�G(�/�L�&�U�J��|���:)y��xHZz�U�ϓB�~<I"V�����Ζ���b�=6��{����)�K�}S�{����4k-��iM`�D}L�'�����03��2����y-Gpq��������%R'΁�5�0��8v�r֗�H\�+���g!��Z���B�u���[�7̼C>�8�sNBn��6���{�z�I��Ơ�lٿ�)F'Sqt�*tS�s��� '�xl�5>$1�@����=�Âl�[I���xo���ݖt�I5�.��٤���l=�0q2��E�T���>�� H��B�߻b�>V��*���Bm�'*��rb�(��ϹU��9l�&͟�e�s���y�ܶH��P ��)>̫ �%���x�x�}���͗�HrzD?ԥ���
3��U��s�E`ǺN�g�eT�,�\6�II�
�:�?Ż	(ޛ������cB��s��
�H\����>#�Kض,� u�棦Ŏ(��|�YZޢK�
ѯ��:?���ٷ�h4)]q~�W�.�x�Q�ݙ����$����ٔ�H�Y��Z�fl��q�k�Vʩ��1���67�巨Mӵ@T_������{��`hP�3�1����3ȣ�����p�C�%C��t�⦋�d�ʹ��S�e[��(���j��O���YoWn��v.b_
���vw��s�^d1���DF5_��6��$��r�IP�jyaP���f����ܑ����uw�b�7��|	ܜ+x����)^#�\"u�l
�ݬ��ͧ��aIZ����)?�!P�P��H�byB*ժ7��/���9�H�:E];�ɊQ��7��a���7�+�R6�V!�C���jw)@��L�P�l�GBL��U[>�C2��ǜ3F��R���赼&�nT},�?g�Kx�->�鰧�Bz�y�U�Ԝ����}j6��E�rQ�����٭��$/n�u�Cv�gC��~���]�¿�]�6i� ���W=ȏI0YQ���zPOD$�Z��Mw�9aaLn�2Ǿz2��eV,z.�>aR���ocۅ���� 
}��A����v�X�\Օ竮�4�5i
�='CP��;�g:�Y�H��E�wZ���Q"�������4����=Ϣ]��@zUo����'^��D�ie��I�� [�^(���û.C�I@ͱ�m�N.]����?�vG������!�o�m(ϳ��z��B��Qb�sԪ�Q
�'�x`w��?Y`��	S\���r�6�}'R��J�g��������m�>^��|d�i{ީ���X���kZ�|)x<�|8h_��y���s�*��K���ǣt�����V�^��t[,i.C�hk�}���Ф�!.�����Z�Ls����XPg	O}*��C�I��Z�F��4�Q��y@l�����z�}7}���h�H�� r������0�1ET�z�j��������+	����
��1���>�H@5P��47;�m�����e�ww6JPa���D{i���뼈�S(�oZXը:qbb����LO	SH�����OEQ�|dw�[�j�����F�+��F�����V��g1�\���9S���Cb�l�"���mR��3�K!��:�A�����9"On����ƍ�m�5�X��H{�9�l��ՕU���Jޙ�N��?!�t:(��l9�8`�o����S*)ֹ�!$��1ca�+ثM+��ཻL�e\��x�����k��hs���w2��-�C�_�M���.��ea��Ƣyݜ�\~^Cx!�>HU#Y4��q?<�{��j���}���df���=�*U#���^�&G���K�vȘ(d��K���F���a�����k����x6?κ��0Xʈ��\������O(�{��`��#�:��,-�9�����+��IU��ģ��QAv�񵏎�txf��(+�|�6��eJ����,��DjKu��c���8��qs ���{]�μGě~����qu~�����B7�4�+�yo�5�"�c��g:?�ů*-E����H:(�)��Uȡ?���O����<@M�����қ��ăҧ�+�|�����L�W�B5_�&��J/��r��b	�x���}lK6�"ުn����	']�e�(-m��>F ���'��.L���I�k�5};��H���B���}����|��ᆬT�ϕ�	�|P��s��*G>��FʎE�D��������&jiw����h})���c���&[U��yD� ��'s��Bk�����S���e��'���<�S��:�ЂB����¶��e)�!hj/�aǦC^ܕ�y��b��qS�V�m����a����F�ӵhғ�\+����A�i��_iAq���6oȨ"S�C��+^���XL��,�?+�y�c��eg�C�)gZ.�17��Ӕ���9m�e��!�YFg�TPNG���5��ϫR�_J[Q��m�$0��p��љ�'DW ��K4���U�7�-��A�- ]������ZX�+�%s�؍oiii��Ï��WY����%X�eH��jS�ڶM*`l�a^�K����v���Z:֛��j����pN�էH���,F�Iצ�`v��F�������*7�L���:��$��lߤ��J��&(̴}~=������sЀ��i߾�D{�d�}�����S�m�����#��vs_8�j{�����p4�v��)0SwcJ{�Hiyy5$�>O���fEUͷ!w3�"��XʴH2�24���3��eiLn�4l4�}� Ԩ�ne��'��c#�#,?�~��XF��&J�)�����NB	�3�����G}29!�f�����wR�|���m�9�-E� rTD��9��G�
�״^��6�G �(�D{��M�p�ƛ�W�G�Z�g@`'�2'?�8G�?5��|�D���ɚ�;	qMA�����hJt�y���k��0���.� ��©B��v�Q�B�̖N�s�&Ƨ@6��T���R�6���y:q�+>�u�����Kq� �� 6㈭{:N���E�|��_۶�&lc�le���կ����7XV[KW���@ ���͒A�9��7����ֵ��8��!�5>��s ���a�6:��l�p47�A`��
����?�^����O-ѵdP@�El_D���tQ/$�pP�*b$�7R0��)��D��l:+����g�2�9y��`��2'��%e�Ę�o߾V����Q�f�4&
zC��Ro��tG��~?ACA�F�a*J�6*�!!g�ܝ·:L�V�QLnJ�ÿN�T��u��b�r����K �G��4��Q�w���{]i�s1�lP�A	�/�����m��F?�s�k�)1ؿ �0��c�9��,��)b�>���2��4��jp���T�U�)�ryc�����X��!�E�c<Q���u&�h`U-��_���~�5�w-y�IS����?�Z����^�};/Hٽ���
�Jݩ5��.��:��h��.>J�C� c��P�6S"��-���4:�Q���j�sʗ��v�0>Oщ:��S�vV:?1n�bB�O����੗#0��Ç Vf�ߎ$�Eu��v�k�����r����z�b(�e�g}`����b��R���Pz�|��!�q$��f� F�� �D�Z��v�y�ׄ� &��:�v����r)h�Q�X�0��Me��2P��
��@��_�C�h����3��R)��V�dӶk��8&�Ο?ъ��]����2�S�����z+�g�W�##�9%��͇���M��Wo �»�(�DT�}�	��ċ�9N�@$F�x^,󜌔�d�P="X/��~�m;� Nd2����a�u9��$/
�����&t>(<��Z��z��؞�g;�Zb�@6�((P���j�p�6�����~�i�F��h���/��*o�0�
7|��ޘ���5kQ`�:�d|O�z3�L�՗V��X�֕$�O���������2YT��F{��F��@��2�j���9��u�~����/3}�����ꍲ�����̭�D�.�e�{e,���J���Lvt+�؁��v�sx"߼f~}C-c��ؘ�������?6�F"�ȳ���8�d��6�����Í�����O5�+p����F`d^����_�xj�lc�D��"H�¶�Cn�z��]����-�?���e�c�g�);rp㜈|��h����8k7&��;�W�_K,��:�¶�~�8�F�t j�h�}��8�������2'��u�O,�����������l��^p	��ے�oi(�j��
��;���Mo�ޠ�tǉ�#w�A���ed�(����
X���rÁP;�*��Z�%�і�y����Ȕ;w� ��=i���B,�*�)j�%]�3#"��ՠ�ۘ�@���W�Z��v��7��g�.#p�ݠ6Bp֔ɡ�[w"­�(���t5���H=�Ｄ#���k�*!y��6��6[�$��"wD G�)�]�0�!�E��� 
(�N�z�6*5�&s5�%�ɇ�萄l��{z8��~�����3{��x��)�z�IY��3bM\�N�9���|/� ��;���0��U0<(��C/ ��ٙ�E��۶1g;�Ԟ$�	��F��6T��m���D%���O�Ű�:0�S��0{���Q] �ҘK�>��L�f��fU��c�p�^�>hX���T�7@}M��=�R���U���xl��۝�j�L�_n��_�)��H(�吻�6c����D�[m���Mz8Pe�� c����t-�M�~8�8�H �vr)�\�����)�1�w����>��Z��32Z/[�=�Z�#�I͞'%ǁ7�w�/t`�� ����a�.R'�ܞ�={/�?�-��#i��+�$�$fG�bD%��0_��*|� ����}|p;�OTu�).�^n��#��%���Lbh�H�GC���{�*Ɍ�{��:�R��4N7���\��#M��Z>�\u���`���"�$�Blh��r�7X� G#
k���uC)Xf��j���t� �����U����.�[�?mB=f��MUd�����E(���P�}ӵ˖���"*���ID�)p��9!�q����g�BTx��W����i�4�2��A��h��4��{�J�����{ԞD(}�Y�F��j|�F)5+��� �ē�� E��������1����]ʖDȊ������JRR��|��6�۱%���*3R�,�c#3���^�w�L<���?}3Z�n&��Ƴ�B�v���e@�6�i2�B'�z[�h��L?ڒ��?%�1�3�}�4qb��t�Sw8R�|ʥC�e>���Z��-�:l���Y���،,C=�����֬uD1��`��{� x�t��ɐ��3�ȇg�&D2��AgR���A&�iԟ�~��B�榪)�I!��gk�%7YА���������rW���˯�Ll!!r��Tk}���="T�Q��۝��Σ5�/�e��_�tK~&W���ݩ28�����Q�:c��mҲ�/��Y�Z�Ny߻�'��5�����e�ꐼ�㆚sũaQ�W"NW��\kk[NG'�̋{E�Q���c��(�sV� -	Hjr])"8P�Լ�=Z�Hgw�OG�}e2�$ء�Υ��+[��Y�˔�!��Oqq���1�J��..��_��=�D��.�:Ku/��o���);O����;QR��oHI9T[�����f���U�N�%Wߠ�?�!	�J�_�h�A�:̬Â<&*��y�X�Y���oU�S�H�6�Z�1��DU�!�)���N{��<f�K���Y��_^(��'D��p���	d8R]K�d�2z��~/\jEΘ1��W�˟��v;v�=�ϼ/#��K�0�S����۾WlyƑ?�K�@�%+�'�WG,�&~H�-����Uo��d<U�wZ�y5p���ߛ����Bh�Tnv/a	F�i�7!�|�Hgț���le�Z���(��KO�]r��xB����_��=پĻ;b#�{�r����b��\��l	l�M�CWBx������l's�<�pV0͍<ބ�,䰬9RZw�"<,FLX뭸�ci��S�K�@��[5p�N����?���k��&���Ѵf��\�7������%�p4Y`�b�Ȑ�����K�xo����4T1��ZQ��4�� ��n�:�6�?�r��H5��9��r�L�}�o���}gn��c��x�?d{���3��-�^C�n�
k�(G��K^��}�`�����}g�4&��AbG7����R6i��ތJ��:�s�����*���C�J��&ࢍ��\�����p'�S����@i>R��H+_DV��x���5�Rêml[H��ٝq58����'�#� �B�\G
�3��qL� ���Hu�6
-��Ƽ��*4�L���Y��2's.�ņ��	�Yu��4>h �3$�hQ�2�|�,�w(��s!�U�a���'g���о�*l�=^�-V8�V�ի̈т����IWo�I�(j� Ch�#��S{�RX��#��T#��/��	� �OL����ؾ�l���G����������v
.�&)�����k8�����OF�iKa���*a�5�6�gTU��2	�B����¶A��ot�J��$��A����a�K:`���h佁7���@ϡF��Y2̚r��*�e�@?��:���"�����mڐ�t��n(���O� L������:*c��;�F+�:���؍���3�RV�O�;8�zo���qd�q���B&�lGp���uM�\��#�f���b-���� �[[���F�c�ć��s��c��Y2B��'O�e�x/n����R׆\�=_� �`��~J�Z,���<�3�ֻ>`,� P��R��� �k=A<7�O���R�%��1���:�9M�By��%�H��j�RqD�&"b���ޙD�:�Q�E>���-���r ���ٳ��o��%0)���z�r�j9e���ͻv��͛8���8����;���S��ڽ��\�7��sqWGG���U�{%�����Do��-���Y�Ŵo���u��t��r
���$ ���E*���n�.Nc�eA��ro^���])1!b��j��aZHyg�+�O����c?zK��l�L�1��%��S��9�$> x�Β���NAN�p_��$�YD��`�n�*�[+��) ~?zN=��� ���k3+P�ų����x_�$���-H,׸c��sZ����!��ٮ�z�Wa`��_N���]�	��=�3'�EU������{�rN8I��਀q�pl�&R��\��,ćuw���Y��W|7݆)�@ٱ��>]�j�S������3Ѓ��_�٭�I�&�U\����{��4'i�:6Bp�u܄,�#ջ�i���hk�]E� ���G���ꁊ��x��5e��Tu�&4�����L?
P _��g+V�HED�=p�Y:��!C�~W��o[���1>���%5�< ����u���z ��3�S���(f5e��?��)�b�_̋��VGlҐ����Z�E5�Gb���2�����N�MK��[vحb�Ӛ���j �^�Z�ߊ8��p����˧a�ὁ��._ظ���Eo��X��X����F�����fu�0V@�m��í@�v�zmԲ�����+b�;�5(���D16��A �9�V�(�	�b��DI�ޥyU��\ԛ�.���}�]�q*SM!T�-?�e���"����2�4>�_ab�;;%�IH:����W�Z=�?s�b��Jcc�Gc����^p���@����ێ��S(�[r�%�:=A�s����m��_�Q��bjܴ���Ks�ki���a��z�_�s�9�gϦ<�h���6�IБ����9ڼM���9��q���ֽ�R�h�wdz���O)�dJ�
���h,��^K^���m���NhJ�v�
N+�^�0�)���c%��%��RI��Z>�6\)�+x�w��yw��@H�n)��Ȱ~&h��G��+��Y�ؘ��+��]f�R���)�[%7��G�W�:��o��*�1�J�H�)������î��Hb�/�Z$�
D�W#�ᢍ&A�+Sb��E0�ٖP��o}7�,SBb����eaD�f?-8��9Xjϼg��D�������������aQu��C#=���� �(�%� �*Hww  !� �Hw	
Jw�twgx����>
g���/�Z�xQ)�f�=�ۧ_��6��Z6�G�u�1��gŚ�Er��5�0�3e`;�G,>��4��&+b:�Oq�s��h�|S���o^#H����Q�2�u�g!��+3�~�M����)���Q��y��������\F�Ǯh����^��Lq�h�u��hL�T!&j��8�>�5w+��䉐��:���.��p���\~,�"B�%��J��A��K1�/Rx���0�JK�X�fXP�A��"�#���V���KO����Q(��*o~k��4�I��վK���/9����z=R8���6q������m���w�rX�
Y�.pZ�;A윢�7�/�ȸ�7❾�a8L�O�#-*�q�R? {e��,����h	���`S���,��C��7Ht�%�{DV�ܐv3+/)��V�I��/��l0��X��>�G����b ����>���Tx�XtTxQ7��x
7��4�]�=5�O�F���ъp����7"F�4Ӄ�Wst1yk&�sj?�ТH���UG��4�L$�C�	���N��;��?ǽ7G�`��c�-�gG�L������ ���b9�5�O��zQ��ʮ�X�{!���Rk��_OU�қ�3-�ۀ���a_XPغ$<�L�m���7~�`r��D���˿Nőbq�9?�:���z��{ؾ1��̌�Fv�Wph���е�1�����@�ֹ��)L�/��w���Gp;I�X��q�\��m��#QL�����~��"� EQ]Okf'����Ӟ��p��9󛵜�,��� �w�3��м�7��s/��ҭ�iAd4��_��_Y�Ϣ�W�Z���A�,�����f@��G'f�v���8���'���@��mL�r�8}�eɸ�F
J�)�!wL�3��lh��FË�tАP���$7���o�{2u���|�D����l]����@11��UC���1Oچ���-Q*��B��pERJ6(��Y��v�%a�3�����V��.�YH���}����Q>�/�����ˎ�J�:�v:��c n}Pw�Q@�2f��!^��֏l�s��3�?����_?�����h��5�3GD�k�v��S�G(~�LY*;����CKm��k4���{`�DK���>����CG���Z�㆞X_�y~�Qͩ��V��!0�����#;⋿����g�LC1I�e�|���w.�iD:�f(W��y�t���*�]i��&<�T�����niJ�[�'U�̻������N��0 L% ��><
WPc(_�˚%�H~���o�ۇ�!.msa�RU��D4w�ԇ�o%�h�͋��k]GU�Qg[1]G��J��яu��f/۞���uH�zN1��x �������(�xd��b׻�z�3��l�2	V���w�-�Y�
{-0CO�F�i^�^ FbF��,}f��-p������⠓[+�Y��/.Ѥ�z>����G#^�	W�L[�sl{C�k��K�;&��^9x2\�K�ĕ*x0�-P�8m�sg�I�6y�je��7�g��`��_Fh��\
#��v���-K��Dr}k#������x�q�b&Q�-]Zx���i���&oV��w��U^��O]��z�$����C����>	��D\������u��O�%XY�f Hw�ij�����62���� �����������Q�  �~��Uqs{���k�69�I��Ȯ�L�9���D��9�>N�2\������,�}�L�K���|Q䋴Q�V�K���g ��״M�Bs�`�G�U�}.5� P�D���d��FG�bN)�Q*dZ��gfW"�o��#E��0��x�#���!
L���~<B��C����@��xz��!ܳݧ��$e;�c���-9���S�9�Z��p�鑦��ߛ�a���Ot�~G��ËhNۖ�",�<λI��!��q�7ȼ��]� �E>�N�����3�Ͼ���vb��K���{�g�	��ꔥ(G%�a�^��m�ppöa;. (�j�u>G�?9��A_en��D��7F��0Z\F9i�l�$�����e�/0��(��AI�h��Z_~~&%����ߛ����w>h��뜂�ɶ�Z���`���|@�GT�|ⓨ�|� �M�x"3�6�HQeΤ�j�bVHjE1<r��g����~�&����@�n�t����%U~q�}��! ���j�2z�I>�K��+3u[n܄?�����2� ��+�M��{kq�n�a{_�t+X�R(��h�CY�#�|�F�[�"�D�3�q2_��9��R��i��P�g��2��l�4���΢�/�x	��]��L��^��j��H�Z�;'��Z�Tre<�?�o:Ԝ<j/��n�Wq��!`-�|/�?ۤ��i����a�m	Dw9:�ȩUu�6�w.eh�Tw���P	]غ�/�&a�߲;�H%{_�f�G��!yqӴp'��wzzL���pE���_T�K��rM�Tl�������F-zp�M��w����V*u����ڧe�Z�7xa%02� ��!��J���D
5���1ey��f4������㮩��moN߹���!o�����W�u�gg�"X#k��B�sl=����Dk�$I��}�6yܪ��=�e7Sad4���a1�~�oȍ��5kAY{᫼�H$Д���(v1b��S8ژ�ʮp$�^"�YOn+3��b�=C�u�����Awͅ�@q��MP|�}�4#�\�=�?C%��7����-+�kCk�KG����#͟m��Y�������P�ͤr�ۼuy�KV��}[��r�q���k� %�UB��C?�"\�Vd��ͷ��#0"�i�=T�z��9_�~؇=�Ć@�$��N�f����PI�@�É O�I B5�7�Z��'��j�0Q1W:�ǹ@ M����پ@�>}C;��2�(O�o*���n#틅��4�o�Lpپu"�fl�7R�6 lq�a���eg�v���C��<C���藥��.�>_4��������0���H��΅ ),�C+�#:7y�v;��_Gt �J���`�/��~��*� {����a7!�t�a8�A䣎�������K F�(�
�#%��W&���O_`�6A|ǫe��tq��.��6�p!�L�>�Ǫ'� �J�#g�o��^ſQ�8��退��v$���3�%|��D�"W��I!����?|%-�5��)������o`�F�q�����v?,�����B j��7�F���<�T?Fk��!&$_t��mޭ�u[" [����׮9���3sb��[��"�oF�C�%��YK��י�7D������!�������ɲv�}�qHVc@üϘ�/��VEG�o���]l{!���j����64j�-��Ͼ=$��;�]��?���\��������`$�2�}�3�[���u2����v�l^!����4�k����P]����O�s�X�r�1����`S����@�oc���`aۤm�f�S�؁����C��pzUd���Ji,���pF�_��%c������f�~w�tJK7L[X�����g����l$U5;sP%xb�������=���M�s�ݴ��q�ge^jkp?9���;��������'�����xDK2� �w.�s�W���ԒQ��yӬn��k��<q���x��c�	<X�J�b7E��]R�Z��P��"Q���'@N��<[��n�>���d��Rq����-d�Eh����+�ᦚ��Ƞ��Պ�Fd�y�
)���Syop����٫�V(5�����>&����rPր��~�x��B�5�Аkg�W�����x�.��
�94y�n�,�u�,c��M��[{����2��������R\�������ƕ���D���K��_N�.�=
8��6���y0��D<n�r9��C�-���u��$�@ej�!|�"��T�)��x�����T���8>g7u���O0�݄W�XAXb]�'NQ�͏f��\��E[NI�׺"h��q���͙�\�*l��B���q;U�#mb��7`�6����V�+�v�ށ�Sg�Y1^��hBE}0wH���\��u�ȸ��,غ�D,A����+��0~M�� ������jݨ�A�Gطտ鏆�p��Hk��6A%���w}���q�U���h����!]̳e��������Lx4�8]�*��ˡ"�b��a�q�*i%�V����P���N�n$,��x�����i�D�٥��S�a��������gk�b��g n�j��<o���i3�5��h�>����W�ŕ��:�#�h[]g��7�Y�w����Ov���bG�j����u+��ڻ�����~���r���mR�o�b���j̪)n}�E�>���5a5>Ӆ��
V2+g^2��)6�N��z�"#`�����%R�<9?0i�WG�2���[�i@��>���ܝ��r��P����p}yǙ�㽣��.ix�G�2���C�@&�^)�~^k���0UkE�G-�8b���/nb�Pk����USC�R�`�gEh�cpe8��U��;�J��A�b$��H`���ǈ��<���[�h��A�F�. �('w|2C/hω�,���q�P��Ȼˮm����YO�h�7�'�\Q��o-�G�Z���vw�
�����8�9����7�8\N��O�z�ic��7Ӿ)�}�F�/���yx�>�A���_7�y6�T�l��f��
*���ց߇+g$$7zK�����M:6�ğ||	��F�*(%���i�j[�Ov4N����Ί�<ќGp�P��=H�U�������*<�?���ono�KH�|��D/\O�NL�=9�sN�Kf���ct՛��k��=�`8	b^���s�6tMuc %2���%��H�_�����P�̩�P���;`n̟en�k�Uod�?�.V�%_��ք��g��=���\L��ɤ���}l�����R�uYpdM��Z:�����.i3���:�vy�}y�Q]��?�g��n!i��D�Ɏ��~�r�ɠ��B���02�r�0���Ǔ`�[��r����L ����j���C���l슲=#i/e7/�[�୦�;���w̰�TS��ð�Sb����R���Ch�R:���#7IWw�M���W7�-��q�5�L�|L�O3^�����L.��_�㞙k��c	gC;�*3�'u�U٢�_���1%�l����h�Zkn1�[��Q�O]���]���ۊ���|��[��4�u���Ǟ0c�##^�i��I:�y&f�Q@"�kQ��70�9�`��t,��#_�a(M��U�4{=��J7b�(#4`���<���,4��<���J�|:��X�Y��̈hFa�9�6	b4%dA} n3L��7SO��.?l�F�{^�5���k�^4�G���R���θ�-���I^�,I��C���v���t):��6̳<�I�����I���fo�V�h��UB�J�4��F��D��h�eS����~gg�7K}�>;9+�&:I,��C���!,{�3���ﰟyzz
���>W|_�5)!9���#|��΃�=�]E[�M��#V��e�s�=��=���`��X_T ũ����Q�����Z�e?��X����3���̶s��T���8�����.�RK}l]M�s�c��k�g�^,�vkK�(��X�f��ȕ�l�3���5]��pY������1{}�ynD�i=�|;��M/��FGҶ8X���С�Fٽ&?���^���c�:ۗ��9͍���&����>�B� j�a:�,�}��Bj�W��Kk�d-�	c�{�A�4���~|�B.��T�-n�	��.gC�I�|.��C�� 3Q&�3��p;��$����#F��/�Ҳ�0�a\^�eeU��ޠǞ��K������r���X�*��P뺠wW{l����km4��R��y�x�琞�X2D EY�y�{k�(�N�O�W(l8�;L�''�jCg��?>5T;����h��С��k��L����xP�j��$�У&������t���ND�(���Mq_N�������F���<h�D8ϲ��X�	:����*^���||�m\���R���]�uvs��(��>�#�;q��/�0_��&_����r=��.��v�U
w����,��.�@����Te�h���y�'�� 4ߦ�3��T�������@�S��3;��$;�$x_27�G2�D^z5ܽ����ߺ���˳e�r{�N�6�
��v�RK�x' ���=87�,�vw��1ߜq9%R���Ǟ�ck{��v>8��٠KYc�ƌ�$x�z����D(��߸Ƅ ��oH����C5��c��E���AՓ�7Q��{�O$f��N+���1n���lg�<6?(O`�S�~�����L��7a%s:j��q}bTON7��϶d����)�a]������F�ߣ$$�`� �ym�$d��ƪ~�9C�l��}1	ni�CQh�Q�<���*g��=�����3���']��S*{8N�0߆&�BH���8����|�����ȿ9�mT��r�U��U�+֨�D><�#z��ͥ�h�i7+���y�#�%� @�[>v��E�T���[i��.��JXp���2������>����k�)Є���Bˆ9�K���#�$:a�%Q���m��H2����r����bN�t8� P2�`��*�[��*�ޥ��X�@
�8r��ԍ�!U��硭�-S# }�t-���a�Y����؄� III怚�Q���&@�oO8���9up��/M6��8���؎v���{b4y�����@"銽��|�����\��o�U�
�r<rL�Kf���3t�N!�ň�Q�?Eĥ����zHv`v�����X �$T���@��s����p*��kO�v��#M
��B����_$��
έ��l]=��I�a��~��Y���E�����p�H����+�>이D]K|�m��Z�ܒ�Sj��)��bi_F��LUUuɾa,R�dc0C����:����S8�b�����쑫��켩C�@} �xw��s�d�tO �7S5����-���)n�T�W�p���x;��v��sO�k7F���n����W(�/�&dj-¶�g��6��h厩�b��F'm�~9���e0ITB�ί�5�Aj}xݲcar����8���U�� =�'�VjtI�@��D�++��C�@��'-���`��W��Y9M�w~��!����w,�ы&���0�w�J˶�&������o����M�U�����BPl��-a�L�d�́���;�X����D����k�t/E�rN|o3����|H��j���.Qb�X&�JW�r��{�	�8�@����.h��v'�b�hP������̅�j}���e/i��	F�Y�˭?�g�^�.M�1��[>���?ӫ?�z�FQ��P�(��9a�ԝ˜$bYTe/-�D���HJ���v�$b.�p|)��:)�J������?L�^�nf�SF��@���M��p� 땆�uqs�"D�$w�0܀�!:#�����潇E-%�I��}c�K��a����;����;J��G�~�\��������a��k2w�� �x�f��Ƨ�"�p����h]c���>�5�?~c8���u��=�M��P1� ���H�B���w*)\;�PG��y��mw�?�����{��Hq�d.�I&�kl���z�]�a�\�l0�gh�34*s����t�#�� �y��<��s(����v =������Y��8������7��#F�a,<���C^�b" K��}������s:[���#����F*֑%���(D
��Zs��F��p���e��f��u(���7��/�����,����R�BH�y(,���)�p�3��8���6`W���F���2[�i�I=�:�(��P؟Ae��<_Z����J�1���R����fm-LݼO�v�O/���?�&�4��R�aB�B�ϻŨ/����'�i�p�P�r����Q�B��RC9:X?}i�E�d4I}�R #�h��ⲅ�y�u�*�bڒ�y7Q9ҩ��b��J�^ڰ��lv3n
�eypPU�	���SUUe���y ##C�C�� ��n^w����ܾ��2~���s'c�[��\��\|C�7::@i� ֕��mI�F�΀�L!7��:UOeF�Y�r���M��Y툺A�]%�F��z�etϞR��0(��am�f<U�s\���*8W���y����Ï�'���W� �;�A���u���j�ߞ�|�.���|�Is�7�'�(�͉����P]uo2#�A~���t*���x��Rm�D��п/4p�ψ:&��K�S������x�=�쥼�-�����dt_�v�~�a}�8_�y5��(���/�{h�c�����d�'�G��M+3F�\gW�A��%���0-B72!�u�47���t�^w��9��My�+uY	���h��1災R�wF����^R`���<��w𼫵V��ܺ�{z��8�˾3v}�H�{���Y3����~�:�<�&6�n* �/5��q��Q�~�4�q�^�F��yG�������&" �^�����6�1�q!���y�����j��p�*"ˊBSK��nv�	(rp�eh6��� t�D��:�QJ+�J�yِ^��p;�^�T;cP[�)��w����A��T7
W#:_���v��{.@�}A�!��	�|����C8F��N
_z�1~&��=�jP)tX��Ŷ[����q;���Gɔq���k(��.�i3\e��Zs��f:���siQ��!�[���QJ�;� ���txے�#�������M��������{5����zk���p��v��� {�k�͑�͠�M�}��Av �8)"��͝��2��C3�B_}#�{���?�&r�8�����?)")y�2]-�����t `+�\*{��^�AN��S�S�?��x=T-��1�Ò-���C�O+~=)E�B*�«<�[�֘N9��^Nd
=Z�i�Y{��`]��s%��T��_|��x�+��+8�-� �==�hbV�dµ�U��e�����.ǗM�,5�i����1��O~P�hx����D�MWF���FȑAH��{�A}a���L�T� [�$h�S�p�	*� �?f��QVT��/�4��q|��7y ��j�#,(P$������?��hm��!���x�$�f����VP����v���u�,�:��?__�N��K�����ma������V`>����Ň@l���x843��M0W`��mJ��@H}f�Վ�l�Y���h4��Sq�:��y����ם9?2�*�@��niZ���@��=�_�ż�s\e�E�yW�=A/���t8�$�SP\ش04��"����8�ϑ@��K���Y��\��� X���������}�X�3B��J�6H����=�l��r�µsۤ�]�41B�$�����
��w&�3�IlםM~޾~{�z�ֆ+l@�Ȳ̆8��'9/��\&K�����u�_+ ��J�)�Y��?�IV��3 �%5?*
�M��W#�?5G��[5-��NFl2�ܻ���r����wC]�ܷ��H.o�&�c�}M�ݟ[���u���+��p���t���CCǐ�zUȅ��݃ǒ ������l�3_I|�K�%����/��[�Fˊ�r^O��!��6�D:P���+��ebĨ��d��Z{�;� �cr#�hy�6݁����(�w��1X�b��(q�����T��ق�˝>J�O�k�;.YC�j�s���I��W�G�Ǭ�[�;��6�r�M �1n@o ��ԅ]Ãw��ԋ�]�oZ<N��X��%�O݅�!�3�A�\���~c5[{G2!��YIA���t	B�RR���!ū�.�$H�F�j��>�v
���˦�"��&��H;�lڥ�'��[�5�c}�pmr>DF�:�j�����^,��Ș�O���<%�L&� ��aA�F��� ߙ�%��寧k��f Q70��v�\Rr��������k� �،�g�-s͐�v���� �S��`���㋐�{����GV弜RĨ�"�1K��J?��k~�~:\�#����Y6YT���(������wd�W�c*�ĸl!�Ғ~@/�u�c���c`��!�Zb�
	�I���I��zy�gi+���T������t���6㈋��̧OY�5���6��fJ�
Y�Pb�8�3�_��zƇ�j������y/�P�a���ir�$hʬ�1��`�#e~*��=e�_k��9�/G��se�/��W3p�󠳗�u�x �I�M��q�F@`��vβ�X��"�{��V��:�ا{�Jz߅0�x�����h沦,S��=�uر�P-V�H�)��J��}m�3ϴ��ǯ��c�d��H�����΂b����������^����~8������Q	k��8��1)���"w��e������J)�f��ss�(�ƤG �?ᾬ�����<�m!�����`���t�zuR���-��Y���/���`�LD�\���.6hy�\5�3���R����鴿���r���U�ap⽷�cg�Yߢ�k��ew��Z�:)0_�3�#F��'5P�+����V�x��A� \WӢYlx�" ��	wvzz��I����S����/�o��J���mY^:>t�I���g�]��-��&iha�r��I$*�MS��g� =�����Ёv��:k��?Q
k�	/F>K6�����Ph����J�����o��/�c��)L�Nv֎� 7�K�n<=oR�(�6�~�dx���ۗ��p��3���%�����1T��P��X[^&#FZ������|�uL�~��y�wo�i��b$u�D���.9>($���v���N��瞂N��|�ʥ�ȇ^>����W)�2I7��FZ�p�S>?B��i��-�EA �ڛ��,����^
]�w)�21r���
�E�e��:O��I����)�_^Է��Q#�3�@? ��4���2�G���~BL'�����g�I_���|�K��'�k3�_�v �M_��'pS�H�����a$����������CIF��H�g��r|ul�W��U\D�WM࿻>���fk�M�"l�_�)���wf�%��J�O��ߒ_�f4�F�IX�ί�b�8��-�Qh ���F>�U��{Sn���Gὃ�_�=o8ͤ&l���H DE[� ��?����S3�t�P���Kp�&�veJ6
�����j�������K~kw� �~��F���d޻�D-�Y_��d���p�L!$߀|��Y����;w���\�l�? �z�F���nc�����[�u���L�c/Ӥ���~����-����u�L�LW4刦�dM��]�іc��O�;���� �H�۞9��}���Gm�]Y��䰏TMq��]�~Q�	q]�ε�+�(��^��k\�Լ y�Hط�YI��d��¨ҩg����[�o1�DGW<�r�a��1�S�{�y������4�6p�<���6$��J����imy��_?NT�)r�/�V�E�>�e���-'e�g����tkKN�F_�n�&����n-�ყ�8�H�`{�D'�=�W
��$�;Λ<�כ�D�R:G�V�>�#5�t6�"�.Y!J���zW��ws���h"�d�εD ����4�k(o���T��%��s)\��K�|��	��znﬖ�f;ț��z�2�ܳerի�F�Dر�6#�Ji��}����j@c��	c�G��M���@��i�ā��r���4��	��<��Rq�F'F+i�ЂO�Zeq%fۋg��#F�`����o���e���y�p�Of.%���x�JC�K�'�ߍ�:���T�0q��<�N�i�p ����l�N:���,�r���b�_\�������%�#��h��KY���4*-==����gc
؃��P�̄�N�W}��#c�+�������8�A��rl@�����L�0�-Ħ�dI�/	�#�S���๥J�,��^w���'	�?�[^y�ΪH&F�������O�L
Ȍ�l��S�iS'M.�"��i�&�nY�Wfi���3a!�R�<��!<P(���dTr��랫��DZ)�,4��u��
0���mݭ�͠��h p�w�w]�6���&Ja�q���"V�"�* ���u ������׬�ͲP:� ��h�q��\���T��gM��-�Z�����Ϡ�����c�=-4 l�u#h�C���6��8����B����JD$�q'ӻ	��!�gO %"�u�>f��~ǂ����,W�9_
 ����t��) ����"SQհt9:�����
��uSI�E�P
9��0_������f�x����D�y�q�B������<Y�SL��#�헢	��ɝ�ˠ;��x	����` �kb�;<��U=#{X�eP�gCd��3Oמꍰ x1/�wqr��Ձ�G=�	�i�Q�h$�'!D��&��4���U؟��:\e�Y��-���N͢B�u�J��w�=LNp̢��!d)��pu!P�u}V>^�N���{?�wf���������&���[=�4��v���݀�׼ծc5[�^�,�y��Z�wlKAwtlA�uII�n�JZ&&��y�̥]m3T����)6:�@o}%���( �$� ���z�G"f�[
0e��E�v�*�ƾ�}���}4{�EV�FN	-P����i��ͯ�'��%��.y�	c
��B���:�_���9لl��#-~O��1|��õ���O�(6�i��E2��u_Nd�ꈤ����v���o.�*�E���o9mc۞�$}hu5r[f:�Q��st�N^�9D��e�;��ߋl��'�`�n
�Qg�)(�z����.U�K~=��@]u�UH��tPO.Ǧ�]r;T$7� h�V)�s翧Z�����Yȅ�ʱ�XlW��_�5_�)O�^���r�ߡ9<Gd>._�����,����K�=VO�j�o" �<�f����
'?[�����@fV��_��L(�`���1n��Du�ev���f��>u�M�K��Ġ��y񫎏��^gJ�bqz�&<��o���^����L���<j{�M�V������B��?�<���i'����y�x$������=�m2��3cw+g�K�%�(�0��.6�kS��:�d�J��b�I7��H�g r�8%
X�*�N��Ԓl8`�8�V�c	�r�q �`j�u��=%����D&(�0jثȱ�����Qw���ad$��wO�HſUi=�s�8"��+QR��ӼF|l�؀��B��,`���/�6�H�;���ph�ٓ�lQ�o��^`�OzF:$� �#�'�p�`������G.<Z-�L����YP-����°5�ⴾ�E��������(�Gɸ�F�+���( �V����x�uf���DD�v�n���&m`�w�b<%~��T�$�&�z[��5>�:�L��.���A�����V�.���ƞp�:F��Bļ�13?<�[�4=�W;CВ��Ӏ���k�M�4�0R���K��R�ה��h[��M�q����I���J-V�o��<�SY��.���9���$�@iSB<�u2$�qtV����a�l���d�TTt=�� <d峛��=��bHW�L��=���t�)��Sz���'�ٖ���,�f��b���,@ڙ�Rư�$��. WjNM9�s֙�a�2^y7����[��\s��6{Qw�
���� �drE�Yf!�df`4D���?��]�l
����ȷo!m����VR��co�`��oeW��o��Vn�
l<,:i�'
a��rM�v�aT�n�0��^��h���ݝ�[o�CtC��?�6�ۓ�PKU���5��Hf�o�(��3�� -�}��>�x���=������%�{J&:���� �Ԋ�q2�_�dzޖWWl�&��D;M^bN�O7��8�U�t������i�f�n��4祉-L��[R�~`І��Dh]��kr���aQ.���y��߷�����ü���~���P
��WB@4|��. �E�CFy���bN��ĥ�^] �}���K&�N���mQ�O�~�y�#@d���+�n�_۾/hmAn�Q=���msI��*�,gk:��ݣ��J���Zd��Y��
J��9M
�o1((	Dq����[k)��>�Knp�jM�C΂�]�6V,�采{��'	��t\�D��g�tEl��H"#K"��wCb�s���нƽ���p� �.���ƨ�D���1�������R�_���ڊU�ڡO����|@�g��#:��q����X�8{�(�~���/�`��&����J�G[��.�3��!��?�3�Oܑ����-��xt��'�]!�'u5�'A�i�v��7�LQNb��$nT\���VDQ��ff�����Qz#������m��+�]��wN�*&mi�ۦ�� 8��%~4(���`_���Ch1���?m�zFN<���*���b�-�`�-�}����Hb�9L�#�`��=��}���Q�F�]D_ɭaJ�Ox�"�L�'���\�{�� #��C���H�,�'�L�ݐR��?@҈���`�����M�"��yΩ�X������d]�Do�ʨ�w�h����U�$�Cp��/�����2�IV�ƚ�箇刧�y�/�� ��W�!�Z������K]���<R!��Qgl��nly��"{��v��=��O^/��Jp.�~k�.'\����q1�?Z�1`����?ͨ�dߪ;�%��?�&�,�f��謁�BG����6�~V���2d^V�pg��,��û�h� |E���Q=�eeŘ�b/|������
�o��ד���jt�ޑ���_��<F0Y�
gy�@
�aq��Cp���?���L>� P��c*dC@_��Bss����;a�'ph�ᢣ���j�����F��9�s�!��7�D�).k����Ɉ�f�)�}�ڌF_�|���1�$�c��-�;�9�l|x:�����u�8[x	���������������¤�s�^�*�!p�s���`^����\��BɌ�R�o�s�)*�=����*}���qK�X�x�0�S�������o<�:+�����1l��!D�s>A~ȇW��މa��Ex�چ����i�w%u�摾Cӥ��Tݫ���?KQ��w��RF�v0	�i��s�јvyS�@]��_���
����G�a�����q�tFP��Z���V��k3t2��_���#���B+��i|u)<��Z�~����I�Q���*��`���������Ⴟ����<� �@��q�߿��R>�{咁.b-�a��t	�Y���I��YdwnY�a���?p�wzXo��#�>k�:3cDV�hy�|�y�2�$�#߅�9R���.p������q��:�d��EǾ��:�ݶ��X��4]#���q6�꫊��g�B	�@Txc�A�j�bb��N630��u�
�efmFEP�A=��>ME~�Xn+��
�#�X��`Y���6��2��S�!��B�����`uK\�tq���;A뛛M�)��l��aM^����o ��p��/�:#�4]3v�pN?I5���_,�`'���+����k̴��K&�}ޅ���[�ݸ���h�ƏЅ�b<.~�֟_��4����_�n VNI���f|&�v�Q��pB�������y3l|,#��Vx�a�< ;kԛo7�F��^�PV������x�o�KF��@
�D[ލ�:7.�|����aQ*ԟZH?��=G1W4#~,��(���3v[t����� �������f���1f����g��'v6���7�Y�-����e���݂x��E.�76-�Ę�X�����a�A�����p�j0��yw`2�\\����o�ٌ�?&�E!3.���` !fV��oP'�Eb��s�b?9e��k_��E9 �X�`��5�5�=;M�޺������	�ŧ1�%Q%�ת%��e���V8�á����T�f��]_(���^U��͈Ȃ����Z]a�n�Ɍ�a����}�61s�&%�ӫUBp�,*�6��^=��n����_���T��JD;�>1��HK�doK�֡���W���h/���a��sL:�4Z8��fa�}���g��ރ��ǐ ���^��x��V^��XG�|����_��aoD���Y��9�bmW��(D����,����_�#�<ߊF��ˣZk�x���G[y+���Z��b��[�EJ6�A���/M]-۴��9Mqu/�=���q�f�`5K[yw[C�a�Lۜ�F��dn �LMQ�(.v��v&��8��� �P�����1z�2`���,�[�).Yc�5p��!::��'#���³F��(��s���j�V��'�4`����^�lpʂn���L�{^�~�ԃw�ӻ�H ��*փ&ip(���*��'��`Ѯ��BH��_)dS�%'ߍ���<�?^��6# %E��Q��lJ��A	%�o_x��|�H�p<�5;j=1Zm��d��g�o^W0
E\BB��-�&/��$xlw[�R!u�AJ];�I�9����zև���o3�]�3sT��t�*°��%���Te�h���y�A ���A(���Vӊ����t��ŵm����̸�Ӫ�j��B;����4����"�N�l����a�Zk���4�gzy$��"ٺ���1�⯽m�SH��ݵVZΚ9��Q�q��k�3�@#eᆰ�JS �@�/�>|�D
C��عЂ��0�4-�X&'Ժ�w�x����L��x^�s��H0aЊj��V���hW^#�EE��BnR�Y����o>u�̆?��~�?��*���H������4H7HJw�t	C�
HHw������%�5�t�����f1K]�zsϹ��Ͻ�=u�.��>C��w�~V�/j�]{	��<_�$x�l)v�����i�Z����vzYwa���Ц�&e:? 3+B:�����<�	��Ӆ8t�s\c�1�B��e�d �w���g�@d���iii�2�3~�|=_���E�1C�x�-�I��}�n�1�m�g�	#$ޛ��/�?0���9��A�����_x&HN ��Jﺉū���ߝ��8V\��~��o1�=����>gZ�0 f^n3JZa5�ʑSN\���)O���\��w�, #k��+�gC�>N��}����v�������B��}cc��A)����O~�uS<D��x]:�TA;P�q���{tP��ǡ)-�Hf?��Ƣ�rd,��%-а���g�5�镕��[� ��n���DL���dҡ�g�6&��_ &1�$�`v��y�"��P[�pf:88؜k�1��$�tƛ����I�QKhC�v?S�J)2�|휷&�SMk��oh�bx����.�"�/����j�ÿ�{�x��~���]�B���ϟ{��Җ�@�R_D��⭤jg3�d-�cJh&�V->iT0�����>y>�i	O[����$����'��Kˡ�`?^ewu�N��-�>�(��		��E)���8�'�w�'G��W\���}v2������L�1��G��3�P�#�^_��Bꌔ����;�v_�o�
L��bo���w��$��(�)�L��87�G���A�~��ߩ�.��B�Q�qq��ݙi\f�SgG\���H9���WKͥ��8���m�hЧ�g|�l�������Y/>q�~NPH��ϟ�dd���o��K_`��=����
�d�c$l��������H����)j@�?�@��x'���vjM���a���e��A:#�����# ��Ĳ!�6 Rt5���W�j�����Y���6%e���K�|ǃ?�QV..��y�ߏ�kl"!d���D�֊U�i�%DoZ#)�k�� eh9v��FR?l��z,�S�DS����&pt&���§��ѥvT��N����=PV2�HC�|��x�X𣖾������Хܢ�ʥ�Nbx�@/ ���UV|U3������暮��l��J+q������i�giW����p_L�[mC�d�3	���3]��I���3�����GYu��N���4�b�<��B�	Ck�j/. I�������G=>r��H��/f��a�ߏ�8@����Z%��O������u�|�_R*�V�4�Z�9�
L�wn�B�\����z��������G����gi��rT"��&�
N)�F��R6�߿�����pVr�!J��//I�L�A��C��

h��@"��q�a���Lir��Y���AN��¶Q���S��ȴ至�=!�f�bV7:����y���U�Z�x�糼״/imM�E*P�CĞ(�v{��CD���W�͓V��(/LVO |��d���tw���)�w-���<�(�
D_xl>O�Q������Pwyϛ(� � �T�/�H�8[)��Oqp�E�>�����a	�}r���3%D��@0�s�C��H|K$d"�����h�r ��<I�¨���@��ǵ�R���()�h��⯃�/��I~�HsGy��T!�2��w\��lI�<^��u3���\Dv��hc+t��Ghz��S�k�~�D��Qe�v+�<c!��T9�O>U�G������Oi ���E��k�J� �@=���X�$�w���=nc�����3<�>_�J��?4y���c��S���/6҃ƭ��ej�(��̗��)��(�7̺9���YR���-ֵ���/^��ϛb�]R<�����4V�'�[2�vyr�W~2y�:���X��((xA���fP9��:�3	��H�����������-F����4F�����U/	�P�P�ʬ6�~zjDѬ,�r-
tG=fZ�!;s��ʇ���T���|���,k�S$Wm�4.WWM�/��ܖ"ccs]Rdp%p�|���J�˨�����#�+}0�� i������Qeɛ~~�����)�c�4"��{��D_g��Q�F����\�%޼�����N&d��j��H�v.��Nb��8y�+19e#��� ��?&�_�l���Ҍ;�<尚���C`Df��q��(���C"~����|��Pރ��ꈣ��`X:�U�y+����ts�Oz���=Z:���U��e���h��N��@!����ϴ��tm?ɘ��n�������kV�\�Ho�����\��U���O�w�/7p�}����
H���U�~w�����PK�� ��=��T�*���2%	���qi���(K��W�p�>V�c��o�Dy�c}�����?�a9�L�u5"w�)�2>��Q����P ���������>�����|\�� �0�G&jj[�8 ZwQ�[3�_3�|��ඕ�p�����m;���?�~#<��HSd{���0�A�Q�!&^��7�b\���^g��Sה��u���l�/ꆾW�ws�t��X���޾/�}N����������M5b Ȑ�ʧ\�{�����>��v�������<��C�.�C��~�q<5^��'+��~�D��S�?���=��@mb���|��#��UIE�)K �s��i�y���x����-qq$�5|F�j4�8F�"v�e>����w���^��(�]r�J(;��8��`h#h<%�r8�s��
��x��9O�K6�L=zɀ�#�����p�1�iwy.�}���X�����7]aV��~��4�D�yOb��#qONv�ȇK��s������TL��P�`zw'�Y9�C:�3 m�0�d@�.� ��<�b�K����J �ܴ�Q��?��3w�ȣ{?���?�E�bO��n��S*�徾Z����I���1l��~Y\.M�0�0`��ϏG�&'�^m;��H�͏h��]����c��Hi/2�\^��9.>^�>����'��,^j�-$��8_�a\�j�2��)�w�O7�~!<��n�/Ȍ����6�O�'����dʖ`��l�����x���o�=.|���2�;z҈Ƴ"h(�3h��:U�J�.��䢚�z(n�NBY\TT��W�gk�G{Y�En���r�5�b�
��N���c��9b�<��o߾M�OSK'�����V_����ż�P�&�}�~��Z*Kf�u��m�qmzs�$SU�����1��0�3
`�Irt�����kx@b?{��`�v�G��G���y�mk4���)k7_�c�nі0��ڒ���<-�~8~iԮd�P�{
��{�N����!;;"�\"��������r�$l<DV;|�TD��F1���K�,��!�E��?sz�I��v}!��O��0�+e�}��S�bi �BN�]�D����p�˷���R/�WLyuόo��*�ՌF��
�>̞7ϴ#Z|Дi�TC9LF�^~9�fu��\�_���g�:�A���ԩ�aBzM{W$��O��{s�/��z��9Z$@Ruĕ�k���U�.^�?�d:g�CLz||<������M�솀O��4t��ͥH3� a�h�/4��m��ɣ&<]~���H�1������N�Ƿh<����f��8c=j�Ак<0��̓O.7�@��ͽ�~d��t7t�#�jJA��J�}V?���b��т�[�����+ș�D{����n�U�F�����J��`���W���X��q]���4L����8�����G���x��ϙg>����A�	���H>��D�Q��f�1����;)i�!!!}��bKj���9 '@�^�~�U��jZݺ�r]i$t��&���gʫ�yfo�F���sKC6D���r������Q��G;ڴ!$�/3^��q?������ͷ��G����+�|��rrr��V���7�B��C�"�@A�7��\����cQp���y���f^��=��}H�2W��շW���9�����+�-FX/���k�R�Ν�L�kq��>�^-�E�Q�����p��Ul@7���fc�L�SP��/)��q%gN�lJ2T?�������Q�oב��Kб4�󦡛�$D�3����
��< ���|���ˤ���l�;&���4S���^���;#�r�)�P����bdJ�'�U���)�rq��Oَ䞒�#�b�~y�E�U[1W;�_�1
����k$�~�R �+�W��>kj�b��j�9�ֽ�i���`��.w�'�E���l��*˳f|�ѽM�|�5�"*���詶��e'��vw��!�i0�G�Ӓ���ދ<+����ـG"�8�4\�S��\o�������?������ȷ��l�`�4��/�*��EY%�30���7h��䮯���7i���K�Ѐ����P�t+6���_�$���7��U���9�F�:�f!Zh������c$U&tW����6��jo;,�T[@��E�z�M�p�J�npa���m�-��]�_'ռ�[N)�Y���͂�B鵵�Nf�y�%Ƨ��OG/�?9���@��£�CC��:�G?��a��P��=�Z��{��#��Z�	�~�S�e���1�Üf9�\L���^E}�a'}���F8E(��{�JTO�Owgj��N��#���<�p/�^�m�������C|��\-�%��̘z���g�z����9�v���/���0�=��h2��~i��E�x=BmZs�y7sTK�sR.Ux� ���λ@��)\A������''a?٣h���|'�z�s��` :�WJ���t�tj�h�l�b�3+�t/)6R�~'ّ��m��O1%2����:V��MI���A��,w�=W�(�"��-Nf���{��{�W���t�1�o׫\�{wއ x8m|F����jr4۞�V5q�K��K����՟�� .5\����7ڟ?��2���h�iRB�%d{���*���`=ս��-� �y�:ۭ�9I���S4�k0	��ѐp�¡|')��e�7�Q!M�&U�>Kt��ԩ��R���������w�l(������лOj�O�kai��j�,t.V�ߖ�n�ۤ��N(=�J��֌�
{;Fܖ�7�OL�:�``�~��P��j	�w��B �����T���#��D>� �d��U"S�&����(����5ճ��.ႍ��ȃA���Ei1e���	0:���rDu���5��O3,��;ekV2�L�|���a@23_��1eТ�? �K�&!��p�L �D�&Iv�����n��-�@`8�%V�X�Y�Xp����Of]G�-�)<�Z�6�k����6Ȑ��.��u2�+�i(M����Ջh�֛���E�b�H����455��h�����[���.'�\��KP�*���@>��tM^��k�BQ�0����,	��P\4���p hf��b���}�v|j�v�#T������ilv:����!ix9?�%���+*7+�~��m|�"_P��ъ�����˭LL��N���e���Ɗ��O�}��k�շ⹸��O0=&�CR���Tt\�mq���I��""E�&*���I��:��E��q7�仇Og�İ��K\�s��
(J�����t+���{��5���+y5���T\0_��I?@F�$|�1����S���I6���H	�G��������Lbͭ���=LL��옹@�e��=k�k�=ufNm���+,w���oOIoN����0w-��a��G�(s����kNJ�i#�%��S��ޫէug=g��� �W�X �>���8Y�� ��
�*|�qT��~\�۪l���|g��&Ilކ@�l���_W�_�#�k�!8�t�O���)�����r���6V��2�dC��K���.yNZ<t�2P�~Vnв�|��3��Ox�3�uZu&�'���9CX2�GJ7`�w���'6��u��&�(�-��=nM]�Z�.������60,�k��++S�߶Vz��2}�\]dh��K�ge7�.�N5� ���G��_��""���|����/T��v�c���3���K�mG�{h��&}n�eo4�x��Ca�Zq�B�~w�Z���x��@�fť��Ѣ��ċ�g���E���&�� 8�$�V��(��䇧�q�Wp�3K,��/�!�vV'N��Y�Ekի����jN���h�q�,��]�`���Q�u�`����]�0����*�&�m]X6�>-��=��t4)����$���C����h�|�����f�{�	������2�Kx�^�	�(�Ά�����V�q)a�'�[i�f��X�45������3�J��H�o��k�!jj����򹫍P�������e��~���P.v5C�2K��>���d,�+cl��A�և{�1� ,a�yۖZ���lcu������r���3l���*��")GYՈ���s���s�A�<^�*���ycRGm�XPe�.�c�A���/)�1#�R�F4�h���85�᛽K4��|�f�(��K������QX�}�r�i��s����R 7� '�[�蹢���^jG�5��UŤ���� #��X�����g��Ѥ
y_FE^M��hW4z���K�z�����l�Ī�T�/M�iR��t�:G_r�Ǻ9G� m�L!l�0j���&��2/�3�g�;|��J��^��D"# ���ʒJ�l��!.�x���d�^�rA�H�%P�#���Gq2��i��G(Ek�U'�Ɖ�*)��G��aE�{Ef�y)�΋��c�G�o�g�DY�$[�?��YǤ����r�������U{3cn�L�$�b`0����IcTɚ��x�U �/�W�p��i�-����������`%��<�:��^�M�l��~�h�G���-�Ǳ�At�G-�������i��רJf����\PT��>t�1����	�o�'''�f�%B����@���>���<uֿsi�RE��&��5T_Ơe��9�Er�𕂆�|�t��$/=�"��d��Ӻqם�̴e��U�c�j��t	4{8������ق?�X���e:K�.h1@��G/������{D`m��k��ĠE�B��Y�ĿC�僗a��H~%/Ai�|��M�O��А���r؁�%�)��z�x�꼷!<9L&�,�2�{�f�&�QJ� \�=	W��9`�}'f�U{9jE��Iys�mc�����3�fkO�= O%#����e;�����IHԓ�ʣpQ��2rA��KJN��h���1IC�nד�K'���4̽���$�\@���c�:M{O���d���?��++Q�/�[I+j7U)t�������|nly�*�1�ݪ�X�ۺ�cmk���IK������\���ã�'���������d�)tI��~D2���@��0T��D���J��fa�yu�BȰP�=�{ �w�C�-�!�gLk�L�
��j�XJ��`���A2y;1.]���,i�N�������7I�;��4O|;�ƷW<Ł�(��*���S�AJE�:;��ڞ8y�$��c�5}�.��@�8������~?��AMW��5ss޽	$a��۫��R��Wi���g�j2��U��4�����Q�WB�Z̈́L��᱌�oX�Ǫ�'�-48�|�"7P�z�S�z�P+����HQQto'F[��?��js�n7�,���W��H/�?�����^m-WC)�E��3H˒dg��f[���)�ٗ}�h�oN����L��?S)%����h�Z�c�3��d�n��T���L@:���HJ(�o�I�Ѹ��Q'66�������-�T=��TI��.%��9��a;��dh��Hl�j��N��e���*Ѝ^.��/�E/ccLt hS2ɷ�C$��_:PE�YҮX���qvP������>����)m<R�E=�0Q�([�Y�!-�+�E���xn�7F��F�����lqx8&���V��ͻ�j��L�[雒�fo�S��wc��
�I��)��F�^{D��A�IF�
�Ý��T%���I]/�`�$x<�Ҹ�M7�0@���R���V��*!��_zD�O͏��z�Ay��cx\PU����϶���D��1���2F��T�a��o'��ֿB~�~�{=�0��5>��)˹n>�.cm�,�Q?U[q�]NU�{.'O�]��j���v!�Z^'#��
�s���G�E����F^Tԓ�������W��MZ{�\+�{F[=C'
X�L�Y���:eí�(6�\]X,����yu���~܍R����^���p��Ԗ46�IdВ���{|�%�n����3�?�l{oO��0�k��t=h�����$3��N�6��V���@,�$��3<{��g��6:���
�cpC���h8�� �v�B��Oڱ��֋��T$loo�jO��`!<�7�? ��o ��yy�Zr��� ^5<�а����vQ��9O��U���?��Pe̙�Kk�2s*>4�j��"��ا�e�BH!��J�p☃ok��G)Y��+��QI��x����Rݸ��i�Ε� 7����M|���MVP�ˮ�x���R�p����O��7)0ӭ�aъ��1:i\�%�Q5����X�^��'3?*W�)BK�T+d��
i�mt�z݈�H�-�������`w��9��]������	�ck�}Џ�o\�$���:���C;ǆ�3����6�'Ono^5��?�J$t���a5%�c�_����q�������3�[N��R��c"55[Z#��ٱuN�a/�t�Б��쩺�S�r�4�ڵ����^蠐/~:�(@���.�?��DDH�ȃJ�Xl4��Y2W��(M�����`��On�a��������4��Ndܯ���c��7SӊG�+�:-�&9��H$�a��5@A�?��RX����8督!�;��I����������DR�5���x?>����_f��/k��6��S#����Y7�wZ��	�%�y���E�g�Q̛�mM���j���ށ�V�C��<3�ga}�����1����*D;{oݴ�����v� y�E�^�Yaal_f#*+��55�k����]�N*2|R�b���u����������=K��i0�H�?7+q_�w���;�B�(�X����NbOrG�xޯlF��j�/�Tf�@�@�VF�Rvo��T��$����J���� ]3ީ֮{j�D�.�Öj� ��^x=Ł���n8w2
��� �HI���D���G�滩Z���G�Ш�m����Sȓ����b��WQO5�	5��x�ܰ��^���s��,y�ge�U���adG�A�e>�ϗ7\�.,"�.��ܯ�D����$��aa#n BJK5x�l�"���%m�p.�p��%�� b�P ��(s�tZڹ]���+Lu��E�sW��7�-2z��ۮ�aV�+�����Z+ZSm����1ԽZ~�M�I@��j�,ΠD���7-ˬxN�k&����m�����}��s��~�\9P���ZZ:����_ŀ���X-�F�V�_F'2<���Kq���O��썞����v��m?ls���d��A�A��<a7�6��u���+�3�k!�E��%��ϸ��j��4)���X-��Q���`�d�t�UR�Y��{���!F/7Fo�j_$]��P��P$[a̬���aU���͔����٦��9ct(	�j�-�9T|�����⽳H��5��t�n�p
��:[��#hY��7���prryik󻼼�I+��`L����F?u��m�V؎�r�����Z��{?9q.�.�zҥ��d'y��^����� ���
���+p@�0��]�=b��D��5f >j,6>��1�j�H��N?�����'�7��Έ������8�"B���S��Y��ۈ�p;Y~��ޑǕZ�����Z�DUT��)R?9dSE�S���@yJ7ʡ���yx�nmd$BIIɎ�ܞ�Wg�|Ǥ��+O��xZ���>��K�穱�ya�wn�q&Рj��Q����ͯ\7���f��0���2|��i�&36#��99��G�Ū�o��ΰ��D��+ʝD�y����#ݖ;�/�h�!��̾)U���f:֤_��p5zH9�j[��q��9���uġ.���Snx�[k�}���SH�n��������/L?L2�ה������5ut/a�q@�\��\b��-�����A(��{�RA�||�_K�
��u�^�������h�EM�HX[�A
"�q$��tsss�@�Wx܋�i�ęёF(�����
M�J�,.|�',����{�M%�S�PeK:�%���\��Ba)�0�w����>԰y�3�ߞ*��vF���%@T��������J���e�Wc�
�!��ā�^z�����1ωT�m�
�qr��bIIԭ�ܲ���b��D�HӬ5����Rͼ7�������ħ�}�.�����)7���n�Xp�b]�i�s�~�e�|Py9�s��%���u��>"a��n쎉)U�M��g���&t�׿���a���6�L�I"��sX�����k�"�����mHaa"FSDx�yKr��9������8}�fI�I�)��.I�2�Io+^|E�t9I��b�ڮ�_���*I#5�����koh�(Ւ���w98�0�3Z-�G�6�v��&Nۀ�{G��?�p��a�N�����&"!����7���0K�{�������5�
Y�r��Ľ��BN;�n���OEXeY#g�m8«��FQk�3�Z��w��2���.6.R]�#�󆊃�+O�E�)��*��i�(���� �ƍ�h��H�o�P�,GU{|�9��^`��Q�X1�S�:S�=�����iF�M��Τ]w�;^����G��Lt����N�檯�k����훧B瞦9Ƈ���L
:��h2��*P��_pZwO�ui���,-�o�b��J�E,�#�.t�w��H;�,&��a�
F!�B��>	�;t�K��R���E����z#�Gc��a���믵CFD ~��]�nԀ�p��i[	�}6a��:)��Xϐ�JR�m��F�tI�G/������Z��5����3�n/����ڳ�|�.5�@�b���y_X��{�:2_̞y7�2�W��������KV��y�D)!�^���{�Ύ}'	~)�د�VbT�gDt�_��}=3��b7lx�S�\����j�x�ڌ�Pz�ډ�"I�r�H h�U����ډ{�P0	(����(������̞t����ЉI�!���W�|�^�bĿ��e;)5�Uj������H��*���w*Ci��5����]��H P�	��#�����\+y咽��-�~l�$i`��$ �p��M�Lڥ�_B�rEb�$�#}8�6�}��,?�x�b�;��[^����\aE��%�Nƫ��OKl�5���$�i�F�����:p��՛l%bԝ�4�@�mE�F[8�(���m���(^��%]�8�AW(w�yN�鈼Ͷ��������#� ��ߙ.� /�����&���aSC����y�dF�<p}9�R���$�,��?�qA��� b&�/���P}���� ��"��)�;k�����R'��.}�n��5����(d�8�
j\Ya�Cn�E~����9�%a�q~M��.�E��+(>���+خ� Jy����k�1EyU:�錶�ؕ��İk���b�N��� ��b�W��7a��b�z��\b`�4Ee��I�c�Uxl���H/+�)�w52?J"Q�J��H̿,u�I�QK���Oqe���r����ם��qiQ~��<�|#�Q��]��i��Hfo<�M���qn
��>�]���4��R��8��mh7z�kP�_b:�W��� ��6G'�b��Y�=v��*��W'��r� :o!/����5��s��k{�>�?� m�o��e���޿4��Ѻ�h���b2�x�,mO�E�W*A��)\�y�9� [�}ND���/���1�y��W%�`�<��?�_:����uC�����=D(IN�� �X.��Z(.x��zL���|��<�I|��(���%���XHk�Q�T�7�٪fs%�������w!F�@�RI��M�q�]��������$�'�F�,�t���{;]���M�t�$k�0��,ѯ*;�@�d�ӵ�4[��9������p]I`���x�8�'�X��"��2�Γ7Ǧ��zM�R����|�
���a�0�m�p)Y��Y�){�<EN��S��Q=��ў_�{���6����*2�=�G��Rzz��m	@xO�s����̀�s�{dO�~x e�_,|ކ�]�t�{�욞��}�A�	�+�.*�P.W)-�[�tZ�
����N��xP[jU0\��SR¨�MUP����諩Nw�Չ�nD���dv���ih �,�a6�+��$���N�p�h�0�Q�_�����|�����T�OFj�kJU0�^��H�Gt����b/U8��R[�4�-�H�r��7� +��>��]�L���;�8�L*D��~CD� 3���?�ȸ�F�R�pn�gۓ$�7�h�����򲸝�$E�}5��R���D���[��~��d����:9���ۉ��+��m����'Ow&'����'8��2g�J��*C23Agi�0��B�),8a>J2�f�M(��km��-^Y��|��v�>gAk���O_�ʶ8N��_9���܊�o慝kx��`.��+.�Ź�svC_�����ݢ�{3-�g;�Y��q��xϦ݅i�7�[��d����F���R��*��R;=j�<	Y"9����ї��Rǣb�hMd{�6���$�`5}'Ǡ��W�@?���#c�>�/g`E�?���W��<�9E�}�[�!���򼤘|���/��dKT��?.Sl�t����Ӗ�;n��q�[��yWT4�{��ypfP�p�^�a�0F���isl(�<��ԩ"�nk �>�4����tu���≄¨�l����	{��B�]��/A6���>���ͪ�xb�%O#YC]�w=e���u��E�˦��\LY�V��f�Z���Gl��V�[��_��Ź�I���y��Z�l�x��DzLԓ��d��e!�{{\t٭��w`���K�1�����.F�wO��kP����72���Pt yL�u�1N�K����}w�iO���.e@�����R˘C*�%��))�a��[_��7y�tn�C�G�]lS&�zZ�B�oO�2��Gy�3,O����팄6j6M��~�����
'>9���I�mpX:�/)�5����	Pܞ�Rw��16e���ZE�)���a���0rܓafL-���R<��v��Tx}oH��d]��`���$���yȁ3켶�^?=��J�B8��wbo��T@1�9��Bv$<�H�h&}�����t�oo�3'g{?f���l�O�	�2�457�s@|>�0��+��^X#������WŰ�:�a7��\�v�3��n��H�A��H>!:!�*��z��� �S��d# ~&�O�|����Ќ�w��
���g��u��Ja5�H���w�r��6�kw5�4������BJ,>uU	/���ߋŦc���<r��R���Y}�C���	M����[�v��Nƀp��uX��̶�<�n7��J��h9����c �&ھ���������V��n�{O�jS҂jQ=�m��t�Y�K��ȁ����-,�����V�]W���Yf�#^v�w�� ���q�y�B�hp���n�����i-�+�㞈>K񅋝 u"��[�.u��a�v?��Y�Vp�͍5���zeT'a6��>���P���B�����������M��/�^��H�w�>#V;�>�{�f��'{�:%�sBÎX ?w��xrs�����:9�����M,Ƹx�.G6cV(fFZ��6Y|O�S�S���WRCY�|��U���[�[L�/��]���f�h���f�${�PZ��7@���p�N���i~��+L�2uQ�M�.�M��ƘXM��*lR��J%y6a��$�BbWV6��;����k~l_( ���f�g�쭞=iK�������\g@=ޜ�>q���!�Q��\<=�\��hlwSm��a?�A�k�p��Vņ��i��C��Y �@c��͇�J����x�X˖��^�_��'^Vų���*�c�ڲ]2]�,/�	޳�r}ߓ6Iy���	���.���;JReгu��ZY��귯��5�7��N�����w]�)�w ץr�Vl,�:�{��y�^F�롽Q���?؜�������cTږ9C;��5�/��Z������m煡��0*�i�Jy8BZ��n�N���xW^/@�H���k���P�[
:���W�\f����!�H�7�<O��o ��7�j��6,��6�J�!Ѝ��>x�wr��N��&0Ө^%���)#֟����
��#R1�w�-�?�֜�q=1��r��)����"�?7����6��d�,������1>g��� ?�T�.�I�\��Y�����46Zk+���R�Ȥ�|��G��5�V��g��I�����c�����L�
��I��l&ڳ��� 0�fI��:z�^�,�{5�H^z���O���e�����b�7ww��*�(���ʂ���۝ �
�����J�6�匢l"���6	�S=���]�%0Cx ��Z���I�� ����^���j�R��cM��xB`B0#^a�^�| N�$Qq���b��gF���l[9��%����t�S׵���~�T�noXP��o�N��
5��lOԓy���o���FE>w��.�v�?����Tn&0Xd�o> ���j}��d �(^�\8q����8�VL}���[ɨ�P.�����j�f�_MbbB������,!�ޘ���x�>��z���a�A2(��ol���y���F�<ŝ���}�; �vW�K�yo�]o�6䭀�U��}���Բ�_�u���*�] ?��\�n�'\�N�HOoT��ao�/��
���ݘ��8M!Ѧ��s���IdK��VBz��1:��F����F�2���'������u���5�w���#��+�V�z�v
6���-�yX����X��z9�L���V�����;|���:	��C�qD��v�r�/7�v��C����X�,������KT]��ug�U�^w��ko 1��3,�����]S�x����V>x��������	F�?�FΌ*�F�p��&~�WS�a��;�+��:�N;J�i#�����`����cީ;�;�Mvׅi.T��8��a)[�3�:��h%�0����O6�՝��9�m���9��j�E��T�Mu9���[K"�0{��NM��ޯ���k����V�_�GR�=/ap��ںw��!�;�~�a9Uܾ@7yO� ��_'��]�Lv��̴��	�4�T�����Ĵ�n!P���3�Rǳ��!������kC�ͥ��f<��/k���1#�+�5%:�`bL0�pߵ�:΄7n-��[��b��|������^�O�4m/:DR��Q��KFΔ�1�}3����9��6�-�`��6n����2H>>��X�^}�P�i߷Wn{Sک[d&��{�!���c���}ia���c7{�R�#v7�e$#Wu��?f�K.0�/n�w$�⫆��x<��\�2��;��מ�Vm�~x�{w��jZ^{��W������
�(�f�"1/�R�M`��ùe�{\;�O�$߇�����vP�3_�dD���]?��w����z�o/�i���Li�o�&=у.�}�xb�����y�VX�Y�T*���Ǌ����s��#6s���qNt�_�Bc��M�8��w�^���v/4�B3�PY�-�u;�Z���{X1x���]
�d�/��׏'<�pq|:c�a�4ɚ��\R��7.������(v��8��Ѝ���~�!N�-�Z����Q�K�ͮ ����Y�3o����N\��M������[->���6X���]�=��;�~��cDOo]Oz7h*��>_h�� ��c�m֌��&]���we�g�V��-$��ŧ��o���>dVYW[ݢ�(�����5�o^�02���u���5_�������]�����&�^$�{˛��;JHtz@�nȮ٦�8q��T����h��֑D,���5,`�8�ݤ :�9�\m��}�m؃�|��1�v��KgO |o��y<��ˠ87�r�݂��).zkõ
N�'&R��J�P����rɉϹ�mq��xz�@��(��!t��&��eR)�&�Q!k�F��t����q�a��Z�(�3�S%�#O�(���B �����O1���*Y��*�UV =����iQ�a㠯,A2z+ŉ�����Y�{�r~º����}"��h�c�gF��i���`t�
q���Uc0��}�d�a���WBBY�UAx�kH�L!Ti7W�J��� �
��x�i�#	�u�Ė���T��7�5́Ar���l$�[j_:zzI�k� �z(��������=e�b/�����s=�x��Tg0�����G(���]b0$Vϴ�m[���s�a�7Qx�%qV>�{' �H����:>�p6�l��Bz#��@6�\��ژ�V���m$RD��2��0��^��2=���:��Ip���������)�vl���@N���y�*BkKf�T��@S��>�		\�+\KuK��J�,j*���ڹ��,�*�bo#O�@�� jB�`���ٱBw�����R��̯�PD~>�i�ax�&���E��Pu���|�
����GU�y�0�Z��1.�<��rD��5��U7��c	�]��!�����ѽr>�\l̮�����y)�ډ{K�5�9}t (��iS!�CG�|��||�Ҭ����;$|��'�۫E���cm��@�H��QF���`��2i��.�iAN�v^�1�S,��:#x-����A���뀇���P�RVv���QFV�we�M����eg��gq��3������{����r�����<�����<��u~�t�;u����ІfB}"���8:j�|�|�Y>PO�2Zg��f�a{u}i����mR�=�
��Eejm�۶�?�����p,p����o.Q�(Z8�c}N�Ͱ�L+�)�Ji1w"-\�HPG�K�ˎ��r�W��T�������CN�y��6PT��k�ED�_&b�l�:��W��4k3j����6�5��3F�>�hT�,"����'��*�Z����Zw��{׼+�*�">߳J/"�]���_�0��\�n΋�ڎ�[�7.����`�'�T�0@߮#<�FR��s+p������pw��.��7�yn�rp�u��o�9��|���`�~K�Ũg#�:?,�~��]���ъnA����W�s�-..��(�:Wf18^�5f����pF�} �h�!0W�Z�N�ga��N-m\���򦪇��Z���v}"H������֓��y�8��Q��e^�D�n�T�,Q�p���^�;x4ڤ������J�����]��+W���:@H��u�u�\N��g��1�!o�RE�r���S>ɼd&ӶZ�ܱ��	;��D}y���f��Х���".��&����P�7�EI7lP3���TM4h|��8�9��kG��	/�DڭNO�d������v�1�{��=:h��|rN��D��s�Uet/b�WY��$�%�)��A꽝ŤI)�Ex�y�_��mJd��Yhʇ�v�d�L0���F����A6U�!�����n��-m��:�?�Mj���x�"��{y)ťqw�'���7�g�>,������_���[�����+o����m�2���mK_C��n:6=ߴ��i��(I�Mb�+�p���X4�o��#
7�m�`���l0k����$�/e�d�^�r��@鴉�V\A�ެ;z��B��V����v�_Y��H��a���+�^7�N����hY�Fq���,���T�_���u

h�K��de���狦S�������j�.\/%��"���J���_��*C�m;���M\�("g��tsi:�H?��q��h<m��=��G@4)�Gn�Xkv��)[D/=^�\~����
�D����m���>�������_�;�%�O�%��sil<e���P?�¦.��ᰞ� �M�ੇ~?�iІ��;}oY�$�3���I.1\&�|�sir��,�I��M��f|�>��GGsu>e|�W�3%˝[�!�6fn�Ա]A�*k�O�_}p�'��@e_�V�zm��<_�����	r��Ĉ�uJ�8 �MB�ZOY�U�ڷ!����Vc�|��O�n�,� �N��nb 2	VV��}��B^^0�}�}w��{'�iLE�iy��4���f�ɇ&�d���2}3��� ^E��(�%%Ϧ4�jK
���Y7��DS��]#!�����r�d��f.ē5��h�~��UH�K9l������AT'�UE�|�}���T&��(-��w����uZW~��3'S:�gi�b�RoWCO���Ȁ�=j/�#�����1 �U/��%����z/��<�$RA�R�����}��%�����U��!Y�sF�����#z_���ݫ+h�\W��q�vsz�A����X��<nwC�Zb#��i�qOf"�+�y��1�<֢\��?F��/e�Pt��5�H��N�h��23��@����	-d"���C���&���o�@R�$-~n��d��o��S���P�4՞|�8ȵ�<�;��tp9ʔ=����C5y���-0"wWñ���2�f�	����VJ�}&���0�%��1A��t�;N�
i2���=\2kR���WI�Jq�|-M�U��ڀ$D�ͳ�1�~�ُ����;n=�-Z�z�r�����g�<H�����������jI:�g���Q�\ˤ7E�.��Tܭl��~��๶U8�+V�{o݄�S�qt�8z����9���d���k�e����y6�o-4wr)S�8�X��������p���ã��ͮ��Ǝe}���>�����{�\�(�M�t��a:;��yW�s!�`��q`��)(�j�G��~O�Ӷ�=pǻ�.���T6nP&�hZYJ}�cr]���Na������¡�fw���Vo���Kz�oڗ������l�:�J}��Xn�����oZ���qˤ�A����|\���h� ��U��Z�S�"��k�������0�!�-.c�BZ���
�i)�9���l��@	>��o�f�{�z�]�߯@N/�&�6�G$6v1ƙ�P��S�`U˫�㔁l\��s��������dM�,���n} ̥���bs���~(R3]22��ɔ�j3g����G�Ϫ�)6�r�S8�
I�L�d����͕�SB�^�����i٩x��@o�+aٽ.�� �L���Yg7j 7}8<���,F��f��lN�a�T�CCxp��B�A͸鐞������j�1D��x�A��B�,�I<�.7U[�jR������qt7�f��o����]fԦ���꠽�)��t^�%�c�7�!a��-]��+ᮮ땏0�c�QoWY�X$�?�1�:e<z����׭S�k�\b��e���i�Q�Inv�ft��o'����Z���|I�mCIo�X��z~�VV�z_zn��g��[�8"HN�_����{E,��D�ߙM^t�Ό6ɸZ�ߐ�E5�DE��d�Qސ�$���H��6�2���X�G�M�e�N��F:j� �x�e��SӈՑ$��󇽿 �tP���)�'R�״��������,^��?S�9Ӱ&��ٞ2���M�;�g�[0ԆTU���|�'�L�	�g\4l:7x�̺֚*�e�v��*�*�v���[����ըK�L-��4m��]-��&�,�o�m�0i�4�|}��(�|�;IDt��� �$���G�]¿�I3��5<hz�������Uӵ��?i�"�z~�Jr�?۩��ZY@�Ѧ*��Ok� �*}� =��D�H�ڄ�E�>��^(g^���u,;s��(S��&K>�qk�2�0~����;!���4!I�<�A���+k}湄� �r��]
�Q�1T�XG\,��SE9gi؀CaWfme��`>C��[Y��F�G�\roy�?y]h�7��ZI��1��a�3<�t��� g��s�� <��Ę8�+��o�G0aWy�y�{���4fc*d�i�|I���z�X��(^$2X/�ei�{a<kX#)��n���ҷ�C����h�؇v"��b�_aB�3R���^$e����G�!*Ė���m ��:5'�u��
 ��U+6���V����_�[�E�	]��%��ds1	�4��Z"����8�h�W>�p�bx~v��6��I&�t�/){���ٞ@t��g�{a�G�,�<cK����Y���A,��&����Q�5*��xے��'�	�IL&�Z�)z2=�5=λ"�<�es�u�H��!P����s�j��E���B��)F4�b5Yl�!�����$�,���M�'Kv�*�m�~�Tr�R�T՗�_�
T^��+���K��fҴk驪	��ЋΦ7��F|�<�IM�����Jpm�����>� �j(j>	�˷�������#�D�����խ���j����/�e�5tBN>%�P�K��E ���䠛[��䆈9�HS�N1�{�.0Z���z����p�b�l1Ҿȶ��/�S�q��sCJ�L["�M�	Ͳ��7�/f��6^�H��,lY�1��8�|��d�a]�n��`�T��o$EN����P^f�^�`m�K��-".�j����.l|3uȷ�?�V�	�N����q�QD��X��)=���`ך���9�����6�VL�����	�j̈́�e���:ʇ�'ׇ��M�x�;��˘_�S�Pq6yi%��n̹�2�L��,x{:D���A0����+��Y��˃���4~}//E������Wc�h;�ʻ�KW*s[	�l��&�`�6	 ���4�C�QC"�zͰ��iz��aIX�uz�C.Qr���A�)�:#��cv�2ī�d�k�C%3ӹ}[AUn����"�k{@�+�m�M-OcA��⁗-ըՊ�.�ayy�>:�Ч�_�tʻaka3�ސ�5�@N�v^t��l��얂b�X�I[0���<E�a �����2߭�:��y|��ɚL���D�s
V�]�J1f�J<��x��O��'�Ϥ&W����C�#BmO�&m���B��5��aBķpJ�,����{��5%%�+��H|��|���|u�M����z�hq�H���`��l�b�FuF�<�,k�����X �*�q��H�Ood	�(U�<as�X�Ѕ×5�`��������ӈ����2�R����zo�����dU��W���|dI��N"k3U6��;����.�;�?�3����j��"6N��q�h���^�E�.�n��g���w{[��դQL���RL����T�V��h� �Օ��:����o�^�h�ɤXeS�z�Ø��Il�T��L�mL5�ɤ)�L6Ӕ3�-G`���qȩ�u8��	b�B����1R�<��!�ݒ<����j
Noz�"9Fĉ�"b:M;�;*��jڴ�
<� �<������ˈ�s����& &]�|u��[�7ӷJ�!YV�� 'U@x5����ՍJ����}q7ǢTGCW��*�Wg��S�}���ȡ���"m�0�";�uX~����|�@ ����ހτ�X�2���ľ�L i��%�4�2����=\P����)f �$�'%;Q��!�n�N]1n�:��y=P�Zd��dNbM�IX���_�~��Q�?���� �|��+ۂ[���cc������Q���==���\����:W��R�w�\v+�"�amnn��⡌׈�6�
�X^]�ڝ�b�p���P��n�BD&�ܾ�H�X�ѱP
G~3�V6��"��j�w��9,\���'E�_5/��ش�9:���b�_�zX�95u��|j��������xR�GA�n�w�Yu�����F|u2�utt2'+��k}�oW���=��} �+�r	)>J	���6a�͍��S�,��O����7���{� �� �����^+�'�����nT*W�8e4CM�ͧ�7D�h@�^	E$�D��t�:-U��č,����}k��^�l����v
$��F�]
�r��?�25�����i/v6d�� /�FútVE�!Ă��w7C����^ݭ<g� k���w�q���ecaL��-���
A�4�ߎ��ë�4GnnXEq}��x��Y,(�J�=n�k��p���e}��Iu���>��ܴ��/�|�������ߍeO5��h��uiB��M ޟ���~��_�DԵe9|Uא
�n��_�n�8Y�<����&0m���s�[e�U�*�"�^sJ*4?;��$���~�- ��o:�bZ�D�ϯ��z�줶WQm�PD�L$F�p�~c�d_{sE~{%������GN��G'��9 �,��,5��񢀧�]�$����=(���A#��j���6��Ze� ���v���nG��s�j��ހ0��[���� �pJ��c|ĸ�컫˪U���y]�EK��D���� �r����:u��r���I֠y��:����RЏNC5�ȇ��.6:@���s��/�V]�B+��C�2�j��Yr~ե�x�S�׼��ܞ'����2�K��Kg��Ov޴LLN�lH5�I53C]�;������	����=����"��w.܀�mjy4�[�dw�Y����2��ɍd�y�(A�=�7bɃt}���x��k9	�f�8]��}���@���������ہ%/�V�2��h�CO�Y���0W��6@�|�n֪�T���W�\9��!A���Ʌ]�^l�ED�?˂j���G {=�(xH'���z&o]�����9���R���3s���kH�Z���!��&�J4�6@����"'D�&%}50�I�s#�:g��_��ؕm���2�E�IQ�+�Mv�-sb�-��A��)A��D�&�Mϯ?z��h�
p�g̟���Yx�d�6�T�"$�xM�m"����E�g^g7��f�� �H��'I�}R��%��4�*���+,��)P����HE��Zc�"���9�`*u	��Ie�kx	��������;ϝF2�,������A4��g?g�@^C~�,�����j�Z�p8_�|�7�;c �۝٢;�����
Gz��
�X��I���?0�:��n'�(� ��Z7oو�mJ��*,0-�ۄX�hz!�7���х���JW�"���q�����F\[(�1MRҕ���h9XrD�j[;�W�v� ��&��o�3A%-7����gʟE��(&$n���O =��d��A�I7$�>��:��I��e���$+%c�C��n��~۩�<A��7�v���߻�b{�NV��3|BÒ�o�vY��_�_��0��	ظ�̃��F=9:Fx��jv��k��`B���c�YTS��Z}��Ao�ވ]�<տ���B{����N��J_ �ַ�`��k�5��>�6���p��0�����f��7�>x���Q�!�3����ϿHE��_��?/�{�]K%����J_��"v>lS��B�e���Y��:>煮p]�0ɉU���l}���GC�u	��ȬL���~-���@\i=�ꊩX;��kd�z����B��lu ������[���T[藒6٨=c|�����N-/;M�ue.`�,+	"!Xtw�<x�ap]:?2 �~��|�j��*�,Ƌ;1
����y��g�)����S7���ZO?+3�y�~�@��,PLKYqP�߹NƉ|�F��!���<���Ɋh=�r����7�Lt�E��Z���.�:����m��:m���^�{�
e��_g|��}�ê�(�E�����|,�-@Ӂi��ܣ鍎`'� M�ZTyr�Zb�q��oї|��|�f^܎��u��&�FĹY5I��ob���wUr�z��B�B�?󏯨�L��
Jf2�_Tde��g�Pv!�od� u��t���0!�F��3F^�=�uAs�*�PgR��j��y���*�X�Z�$c>#�E<l8)��A�ͧ�v��.<�ɝwG����E'����n���Fw2	�5-W�< ��]�jcz���+2��_ޟ y��'���{����Q��]}�����srQ��>��/h�E��ድ��66.���i�&vq#�[Zu%r�D�]�ϐ���0��
�	�5�G�o]Մu��C���o�1c�8�����o�������WO>�v��.�k���T?���%�(2r	]���6�� &-�� '.ϤP���{`�Jjȕ�b�}2�c�������l¨�_b6ڧ�N}I���k�A[��'�_��rn��:�bt�h�N62��W�v]z� S>���A�<�a�^ƭ[b�D����<F��/r���at<F����B+(E�o�x4{\�RcI��a�������Q�SH7yt��=�TB���*���U(O���Z�0�9M2��3�j"v��h=j�ׇ��ߴ ����w�����u�w� }�$�<^�@"+Ѭ��{���K� gR��hI	���R����/����k�~�N�H6�>p��0�` ��ꂰ�Sٺ��4pP�k�K�
|ư��
/������>?
��)���V�=�4@�?��S��L��`�GJ�/s��� ՗�\��x�/Ж��3Ҩ�t׭3V@H=�e�3~����6�:�q��s'tۣA�xp�1�-���3��0P+ZY4�F;�(�n&��U��Ic�ܝ)�Pjz��MO��&��G���σ7���:o6`�X'�6�dcC����J��(�O�,�K�����F�71P��'%u�R�q@�5�"�.��|O-����R�n�����)Qx�{Z�6d��?V���.l��)BY�L���*��`��t�e�z(�]sB`O:K�7V��zkx���{_��[PQ�M��ݡ�b�쉽r��*
 } �J�S˳޲#`rA\�G�+�1����0@������w�8���T��g�+j�!�ċ�b��w�`<��w������l��X H�>��c4ޝ���#(�y�}�:�ȕ&>�F�#J���^�� �i2���@CE�c�Sn!M����Vw�p{~�0s�T[[;<4���F�������c�����*)i����^�a�9�&��?��4̓2�_ޙ�>횏�+9��ϩ��I�q���T�5*]f���t���xFރ�y͉N�|�=���w�y}��gw��n���:Lr+���W}��Mڸ���|Pe;�)4�n3Z�)'���T7Es�՛,�Ҥ���C���4���R��������:4]LyyD��v �"E�/~o��F`�>��f��_\��g�LB>�R�֦� "�wV�?�3�>�9�Y�:�=�^o�dhB������VC��]�%ÙOBL+w��@��*g�qxa  >l��X���M��� rv5E���HH�J��������)���UΓ�� ߓ������_��JgĦ���oN4��=}���u���K� ����g��?^�$�[ 2>@�NJ3���og.^���돹3!�R���{̹�/�.  �A�����&��4�;���m��u[��6#�
���[����\������0Y�1@�{��s ��ЭɷNY�C/�7*f��mΰo&+���"��j08��(cc���䐜_�������"M�kr���)֬{�/%L9��ݐ��3����U90/����S��*�nk�ذ]���V�m��WnH�"5�Y��O�IgyJ �A,4S]u���B
�4�2Fgf{U��5��y4t(�7_�P��V����|_d�V�����Йb��-�i%�����S�#�����8*O�#����򪱞�֛��ȿ���	�s��&�Q
Q9� �T�׾Tl!r��p�Ԉ���Bt�{q+��;���KL����� z+�Da��ޜ♘	P��q�%5~��{���3�D��H#��&U�\�`}������J#���տ��=�
�Q��p�GG�]�\�B��e��(z�PjF&Rc��Ɲ����z� ��=/���~��$2�Q(��U�H@/x1wE��w�,��;0�:��a��m���+���v~�%��i1����B���j`ABҹ���W�Q��<`N�ߙהK?��=�� {I}���Ή�66(;����ˎ�9\yH�)��h7����@s��B9�W5g��ay�b�}`�O�=e�Tq���( �Hc���kH+K`V���H�P(��#%�%�'Pu���T�2��K���m��@��hk��B�͕�����)�c��Z���O�D��������PD4�{

�5� �W4�B��w�R��TӰ8@��nh���\�-�h>0���禽}��.��7N���P�b��L�$�D�ܣ����'��d��S�-�e���� Xm��wC�|�4ђ��M�����H^�hDˇ.����ؖ
�J&�8J��{Iq�r$�5A�`e���*���/��吅w�%��Ǔ\^��O��ho�):1�x�a���/+�	 ��x�]���7�+����c����uL��0�����K��	���q:��_Wצ0WU{ӊvh�w���/P�A�#����K��\�wk��'��B-���>D]~;�{M7��V#U؉�Lj��U�i����z����րr���b~u�Z&���a���zQ��)��Zq���S6�	��e�4��@.b�:�÷��$�EKPQ����#l�q"��՟��.�2���Ф��d8�OkW������U@���o�o��>�>U��_?{�C��b��Z7���::c��R<��2��;�UX�p�����,@����w̝�ô2�����Ƽ^����i.�V��;��������+�ֵR�y��1��5�8)�&��6�|{"�7a2q�e5����t�1���o���@��ؒn��67�%���[b_QQ����Ң��@_�JA ��߽A����<c�t0 Ib��K�p������p+}�W\��ւ��ꟺ��4�m�w'�v	�x���9I9l�T�&�wq�?C�^	Z=o��Ki��=/�:��TPO���^^�W&kA�-F�2�� d!h��4�*7M���=r���(�Th0�jhD��M��<�Ty�Y�
�i�N��6�"y {�FR��p�`A�Sɛ�+vR_{�Y����ɗYu$�EP;�yOFU-wr�T�Ze�`I��NR4��>�Lu@J����U���W�������KH�F����x��ă�#F6^oes��s�!	��a�
U#��� ��o"q���P{y�ԈA~�l�c�U�Xb���|ʵ��P�"ؖ�%�IUR�?	my���?�M]�z.1����m�&�~��p .r�����~��LyL���S=F棗p�OΜ�d#$����KIs��{��\46h*��|8776�|��m���݊�&S��=��6]&��0�����6'�x=�$�d)�j�ޔ��v�lj�]E^Ѝ���\�PU��A�,����uPl����������z��sb��9�k�\�:������Nս�0I�^����ee�Gq����j�Ca���h. %��l6����S���x��-�e\Q]�����>Q�+�?E+�D��x'_V���zM'^c��՟ȑ&�l��������xJL�.	4�nw`�v�;����{�}"�eY9�g�؆g���H��@me�<�v�d�b�oߴ�9��-��I2u�]$9�T��R[�*��Ңw�!�D+G��8s!1A�$���^�^��̛l��j��1�J{F�~�E�M��O�D��D
�����O}1o���g�L6'<�9�J�n�V�M��'�z��<������59�F*���tn�ȆHf���פ	�Mʈb��9��6��
"}U'����C��^��:�����|@A:X����?��8�_cwv �Q�;��>�����%�q2�W�l\U8}���;U���We���,�)IO"z�7#7|��B�rR�$��H5�gT8�5L� �E����k�Z^��k��i�����
ޥL�(0ص���^�V@���ֆ����{i��^�~�v��^���O��
!�v�P$>�u(��Qu���Q�T7"�qj_����4�Go@m0�}�jQg��I1��Ba�eoku�wǦ�[B�����A�SJ
���K���)Il�$�8�����vz�^W�;/W߬p���`{�uó�E�Ed�F�2� ��s�7N�/�|�}����:^�N��!9�j�C=�@8^D]�y黺��Z�3�h��U�I�UKP��^� ze'�(=���p_��Y�(������V����	����8�%/�A�W��ZHA��D����i>�z
���˵� pL?͈��I���*���V���
������m��앁Z��9���bCګ|�)H-Qph�_���-�>�/'�_!#	�?�>��
��Ku�L�a�1.}�?V�?��V�.w�6}�
}le�7���u���Z�H���v�����*������s�Z#$�`M��.y��)��Pq̯B&�4�mH���̝��Oe՟��q�hd�1�W���
�S���;l9�����ߩ�qO}��/E0������(M%��$����5��
���GϢ���;��8�r����w^-���7n�����EV=ͳN�:u�4Sσ��Sg?��X����ts%�We95��#��T����p~f٩�#����9� B��;��'��k6Е��������FzZ�B��Qp=�}D6j\7nz"ԗxW�'� ��B�ȡ@�wd�~=ٲ�5�,{>>ƭB���J�[��fT�������09C?`:�#��މܫ�� _��</I&9������#o�-3����� �913�8��:�S����gz�d��'��/+��IL�Kv�c�N-S��߻Wk��`�Td�sYцg�s$�5�4ԫ઺�_�g}ŧ�n�P]�I�8NW�ꘝ��o?)��[?�}�W_� Q[�9�c�*u��X��㽶
E����������ɃU9n���۟��c�@��������3�)wпﲠ|�v9�Z���.W��Z�fW�l��0���Ɏ��z3�jsyp/�,y��u�Zu-�0��X��4u���m]/*IW�E���:ٖ�s7��-�n3ק��{���c�������Uy��xo�mPR��DFT�!1���F_'YH��.h�������=�.�CZ�<Mx2C����6r�P�#[I=;eǥ��<	!���������?;��멌��WB�y9I���}A�(�ߥd��\H^(|Wl�`���.���\�&B�~�k~�?�и���jY���m�!�-ۈ����5�&���q��Q8.IN�ގ�ȸ�^)Y�	mt��LUW�����.���@�V{}�p�zC/{�ۻmHz�*ِ���c��T���hB�N�x6��^��BfA�5\���_�L;�ÿ��'I�pLwԡ	��sx� ߓ�Wx�Ȩ�U�f�����9�9��J�.�|�=g�rs�4_z$3	6d�c�(Ŝ�>�ۥ3����Q�N�����Tw<'�׭_2�#M�qԼ�޿��%ɒ�D�e��&+�:�\Y.��J)��bn(g�E���D����S������=T<��:]]=����q�Yz�6;���� ��?��`��]q��q�,j:
�l}�J�`;�N�[y����. |�y yD�0Jm���$3}������)�(m��������#��b����ŭ�ٵ7�v\VT���$����j*)Qϗ��|J;�;��U�.{h7�9��a^��g�ŕ�|h�:Y�D��L��9�?�� \�R��=���~&y�qn3.�*_���~��_ě�1��T���V[?i���S�A@ƿo1/M|�b��|�w�H�L���'^��xb~��Բ���|�� �Z_w��6j!���;	����~?Wzד5q�`��æb=�۷N��Uȁ�b}����hϻ�Ѭ�j�-� ��/�<��� �*�P�z�*�撜�S!~n��z;1r����
��j�G
u�8$U�	�F�Y )-��lH���!&���љ��8u��'��9�	-��d�l��]S�n�(����䉇�@r/_ro�^_���EI�NBz�����2��K���hSG���]_���<,܊9{�Ɵ��(�d�pp�3vJ��A�m��q@þ!��ɾf�y�3���c����.�� ��i��[q��)d+掬�N��5���Y�<�<n�����h���.P���Hen�k��aٯo���4�z"�c�,b{:O�ba�om��ƫ@����ǰ@��s(��y��&4�.␋>�ڼ�=!��z`(�i̬�V��t�@y��\4�IDg�jmn��=DA��o�]m�D�.}� JY������`��޴����ë�f>��O�&����C/Q|�{�>�} pc+����5{l���Q���g~3J�C{Txy��l��]��o�w
v5C�n/dx�?6h�2��"]��8��:뿦s7�6Q���P\v�S�����L�h��%z
�l��g"-a��-]��;vNx(�gLB��^�./���Z�8�kێ���D���Sa6������SOo�6�l��<�?a�X�7=Wۃf�C��z��-�JG��n�����>�W5��U�W�P*x9\y�钜s�Xy G���Q�6���^���CM��$`�۲�pԒX~���N�5����I����*A�vA���*uui��<�M /��F �´Aٹ�S,CU�g��쒢7�z��ߊ���e��l&r:KK�X�;>�r���'>!�@�	T�E����5�j�6A|7�Į�����<� }|�<p�{a�t&�*�((�6�ȸ�vsj�G�1hf&$wÃ`4?�?����&��9*88!_�NY�)Q��ѵo�?'�Ky)��aL����⢿�h6���"�'��̒���;�(��+��:�����C��Aw��,��>��X�x��\<ނ�_�oxX;W�i&�j�N���87�w�v��M�I��ů(;yV�m7 ad�+I�<���nr2/�J��Wd�g;&m��f��7p��뚰i�9��B������y�>�cֿv��aW"@��{ٞ����O��E�U&F�QL��������E�n����W�1]Fv��U_���}ŖdB����(�����
)N�x�Ͱ��ޞ?1�8υ����w4�Vve~����#*�,����ObO��,�4W��@�i��CEjZn:mC2��]^]�amD�ܶ^��6$c3}�/��)�z�J��V�0� �Ju�7�>t4/N�6��G�U�Xt�_ /�J�
�'�y
	6yt �>���b�t�<C�T!��y7��ۡ���Mu���4^ݾ"*V��;������2�?����>u�W~$ғbƻ��_z�ۀ�7b����.��N��:���㥜�>�����!~9����bOM�K3cLӁ �G�KV+s[�NZ��5������ʆ�:z��pq�Gb@�����ym�ξ�;�2� �H��FZ�K���c_V�)P5�/oZ��V���&D~_��A�_�K�q���������I�}����C��}�_�>CH�b�M=-c����ybsUI���)�G�lډ�@oW� MH���G�7��`p�d�XQ{A�;F���N>Oc��_ԛH��Ҟ��Ǡ�����T�*4Kq:�o ��aY�;�͕���Ǣ�v/�i }N�,,e�/��_�EG���eU�����$�$����,���C����ي	:_X�@yo��OΫ'��b�i��᱋˫��ڧ6Zԛ)�jwL�?�Hh���~���o�p�Y����
��A
E�.z�״��/�J�=[���,��&)Q��i�:�`lN�|UsE��1%U��r��y��zZB�%��"N�?�,cOy~��a�z���8FOzd� &��Y ��V��T�ݹ�B��($��B,�A}r��&2��t�*��@�%e��Y�sv�q�#�L`�u�<�������1l6�Ŝw݄�ij����7'��I�`���<����2�Yt#��X VY��r=au�:�5:{���tJ.�Ĳ�[����+`6#Ɂ:�]L<sN��`r˜�������� }�x��y�b��%�V^y^� �I�tK&��k{r�`���Oe�=�I�q�j�xbxC4̊��QS��!�=7	�tI�_i��淙&l��s���Y�#0�_�C1@���
�ZRYi�N:�Z �m���b1>Ssl��}��7 j���L�e�Ȣ���<��T���n@�t�|ۖ��e��(���GB�㷾A���~	��~&/eu�p��n���>�,�XZ0��1�'I\��ݵ�L�����y͉ʦ���zy�gq�P��O��=5�1���nCsu$_�S,�xys�뛂t������x\�:���Bi�{fb�Y����B�Ǝ}���Z�?W�'E�7����`a����I���֐{�e^�;�)�R;�1`�4�����,4�L���Y�; y�-9��H@�d\@�
���C�,�:����g��A~���sȶ����4sf�	�����6
��P���P�[��6�p���*_��}� �LN��r�E7��Q�z�5�4C-⸵�\Xa��2ry�(3��!��l3����ex����Y��E��
�s3	`��K���̳|9�������@���IԾ�=е3$i�w^x�����	_���k �h��3�~"����w�'�i�d�vT@�r��G�td�P���B7/�=��������F����5��!,:��E�L�C����ē���^���!z��Z%nƎ�ĥ�7o=ۧ2���t�"}���]��D~~O0M����F�[�=�����iD�q};Ł��>?�{�Wq�+�Za�`��R�.�L���t��s�|C'i~���!GG���F/H��ϖ!��e���.nF����r�nJ�R�4��Z��D��SԔ��Ѹ��t"��@��`����SQbS��o8L���{à��lQh���r�є�����_44F��x�uL�>����X�ȝRl��F��JM�)-:��v`icm��w����L𔯎�ஂKQ�{ko�T8!N�9Y��\a��`�m�4�~vt��C���c�'���N2���e����J�XQs��s�m��綾�h�o������|~�{��rep��dS!m�Ӿ������&j��ӎ��A�]��V (�������=n�41#�R��֨����T�+lv��"k�n���.0zˎ��CV�����E�@dιf������;�:�<���G�G�����/ɏ.Q�*<�1 Y_(�?�؜~6�/�s��?~�Z2��Y/R�P����""�;�F�r#�eh����������JFvWiH���)wZv�kԃp#�a�Â�KZ
�Z0��ʲ����ܧBoL� �4EC�5e��#����	����c|�y�:�8�}���f(��;퇦F�t2��8����_H�V5�/"�j�,�S��2�-x���~��8�<z>�K����J1y����S$�y�&�'��N�8�~ܲk`��_�iU<#�@��2W��ի�8DD�d��I_�'䳶�K���z5��v�a,�CKTZ̏Tɓ�+]J�c���4;���K����k�=�}�HC[7U�@|W�~S���dw�r{z��i$kdRJO�>}nn�kv����>�$�s:��8lv7Ο3�n��E�+s8x�ss�'�Z�x��;���s���X�ܶ�����	ӱn<'�FV�(3ꮪ)K-?�?����{�w�.��)�o쁻�h���lP����Uw�q�P9�ߔ}�_Iz�JcD�
���O��I�/�����^���]��3�"�cD�(�6�ΩgO��Y��@� ư��ho��zS�%���ͲQ�rgC�1ȡ�:�M$	;�3�wI����$#����|����),䀘��V+>��{�D}P�a��	�Gy�7|-�դ(��Ň�bM�˭\0#����
�������

�J)  "��Rҝ"�]K�RJwH�t,"�K�J��Ĳ��]����G�ϽwΜx�{f���BZ�l��t�𣒘>λ�/l7�����-�p��E�`K_S�C-"jW"�"�}���}m���F-!`�2�(Ke�m�*ل�8N|#x��H�Ͽo�����8�m�G"#�{j�F>�w��J�K�L (%��NWD�*��"���s�*�����v�.����b�B��.P�o�w�ٍ��洯�2|�fۀ��O�t�h%
F�ڸ�{���(�1Rf��OM�VܵT&�����s�-���*?�9ُmiiR�9�EJ6�d�6.�����흯�*��F/����C��Z?,wM}	6��e
�Y,{{�c��C����%(�!�I�j��a��Z�|1PG=P���K�z{��p2�'�4Y�pG�5z�{��\O�>���hV7��T�a#�B�*2�����|'M�+á7�J"oh���<d_i��ĸC���8B�
k9�u-��;ic�H:#DS�v	�4�@=��w���N�y��iZ����Oko3�S�/ݳ46�sݒP:z��O;�x���?�|B9άnE%��y{8}n�x�1�O�+#@է7�_���ɭ���c۲*k��)\Y#>%^�
��	
�E����>�=������Gh�]55�\�C�*�]��Ǩ;�&J`_Q1��//޿��y9l~�,� ׽�!"I9S�Cy��+$R���Z6V�/�LUI%�B^�A��S�U2d�������9$�L.%RS�qog��hfz��:�d�;/��Ol\�[.U@��Y���|fC�^�cn����?��t�Y���e7���z���'1z��Νy�M�8�Ɛ�fb��;�֬�m�n��@�(d������q�� ��7V��1�Fj�5�ȅU�����T/��~���ݮ"Y��E��%hK�e?Y���a~7�)���]�_��K���ܿ�6v�G��^'G�7���ל/
%k����o�^l�7~:��۶�K��9`l,j��i�lT�F�����.n�di�@D�7�o��I?V��/.Z|Rl
]
�	̊t9�rg����#��Q�gl����˲�],���A?�EC�s���*N���_s��0�I�!U]C �`���
y���������5�������q���|V���ޛp�����b����@����6���1sT�@�P�a�����$��ϱo�I���=(���!�g�,���$Gj ��S{|_ĳ|É��Q �P��4;��w����$
�K;,ܻ�  1��F܊�MgO�X��h/>�����TmeeK�k��������=w.T%8�P��[g�_�!.�|l5ֿܜy���~�JpmťoϜir��$ w�%N����r��뺞k�,u$Qd�2�]�)�q��B����}�q/�Ǳ�*���_�V�)`E�\k\�Mo�~p{i���g ]�+@��@�Pq �H��VF*���Y�DO�E06Y�<���R7x���~�Ɲ��:_��y�ӡ����+��ݕ��-�/�@�T��W��@Y6�>�Ѳ� I�F� Ni*]s]��E4�笌�M\_7��}nHj\���_썵�U-9iV�V8�h���ml��Z�X�%𖥉��<Fba�B���0�0��Β��+���r�"�r�4�7��OOZBSd��!2�^ֶ4��2�U���Y/��Td�M�~סW�+#�<�U~��AÁA�����:��g�`wE����:a�ruu�Y�Y�@�GF���U�����ڪڏ{��H{�rf���y޾Wk�aý�v�me��qҢ��H�;�	�q�n9��SK�N���s���O Ns������#��V��S����3і��hY�t��F���� ��-�g]�����;���Z������L��Ӷ{�NZ"QJ�����a;d�Fg�X�`]l���5�_Ym!��E���/+�m����ǈ��77+���b:	����^X�p�n�g�m�s=���p~i�vs�K^i��9k��'d4�$�Gc��e��W��h���F�S��&1l�-��*	�	ʴ����R��S�v~��X�(k��2Έ��\�1���d�t����l���fR;du��5q#K8H_P��s�KM��yILa��"e��76L�ǅ��å*Me	P�{/B��J8OG�J`��F�@7$��$�|9���.B�I�i���e%����� �Fy�<3� ;}Eva����Ԍ��ꎗ���V����y+��ݿ~Ud���DЌiG��ގ�OԿTÅ��<��[��z�����":�;"���h��U�!qM]^E�0:p̨����;��[��E�Fl[��"��b^� �ޓq�`P���r@Ho�r���?�򱢿�]�#+CD�!jlFZ,����_;A�o�:�qzX����dH�}��^���_�\��8� �A�*�$hp.PJ�����}�L6��|�<((���%�S������}�SN+JM�U���j���ё!��{���∩Kd����$��ւ�����ۼB����Ȥ�����ew��W\i��FX�<l=@��1��ep��d�
b��cG-�x0n��&���f��	��Z������X�� �G0>�5谎6&�4�xa�H�2���>�=���-pGhdH���B��d!��ƕ9�N�����8z=��eP�����j���kmS]�=�?������E�'=�F9ؤ��W��4�d�HZv(�>��T���^������B�ߟ~�\-�>��rtu�����9b*=b�d��э��@U칧Ģ|��s�4���s{~��/ɭT~T�^'�����-P�� �x�6���w�.�񗞽)p�PJ�������E%��NQcR��ٲey�઱h^K	�a]?æ�3��]2��X1��Nr��Ip�����G��ŏ�"E��>"�NH��'h�,�r�-p���/^Rɽ���W�*�a��t=vrxX��$63S�:���o����T{m�q�
�nU�Dda�n�ݱռŦ��X���奘���T�?��x\O��a�BT��$ڛ��=�?=�3��%ɋ[��-�*��cqɍ] ��_*�������؉����h��w�H6��]�04S~�T�m�>d�
em~G���.��T��:'����A�Df�w8�=�� ����XD��5��Wz��Y��)qNꪕ��plo���٬�Wu��c�=j�}�����D��t zNj�~�I��d�z�.	H� �qtY�N8���'6-�tu����s�z����^�����8�`ä���>m@�ԉB��*S�죏^�S��]��i�0}5�X�;���	�|��+mm��2W��F�����H�8���I�?fb��$�A^#������++U3�E=�fk_s���I�9�����@�I3C�E�$%��a�h���$�B��!������;�V�����rC��U�W�J��ӧ�n�/��T>�0,���{R��Wdm�0�v��ѳ��b\{�����jp�S�n�� �H���@D7�{��6R�|��(��kW��G����e�I�n���"��� �,,,윜J]]]����yx׻��ʍ�r�Y�]:�I�3�](�.��+~��t�23(X�C�9)ثGT�a<��%��1T�!�XK��(y�R��wxv ��������YE��4����Gt)�m�_��^e'�^�K�(�V5��&�j����Z3#�kI��WvI���8F6;�����9���&�$�t1�ȏ	]��]��.�u���46.�ܝ��=P���I��"CB.99I$[��y�7E�0�r{ccF�k5��m�ׇA�[D@%s��Xp�o�kAxr���&���fk�qI1l�hp'��o�0
�$�/�� ���-55��@\�fj�`V�p+ qZ�����i�9��Ь9G��ԬS�Z�<FG
}(ε
��]�5f�ݗ��}�?�x�c�`f{N��"�v��17������ϼ����W6����E?~xݹ�����0�B���T�j�G���*=����Dp�Yw�u����,�A<|��<�9�4��� ��e���y)�snlP0��a�<n�ee��_0G�
(�4�"�D�v9�A���a:)%PdJ��?�xr$�^5��4�3U0�tW�4Q���ʩ`�
B�8�?9�k��As7����Hr����������	��2�Ce12�$p@���]O[ ��W΄�*����Ǉ�( �~W�����Ғ�Ȧ�t�X�6W��?�
�k� L���ș�"����U ����y�M㎏�7��9�
��_�57(��f>ޛ��\Ҩz`�A�g������*���'>n�p$>:%����j����k{��^�������gc�/ƍ��zl���z����"xm��@�(��7�OOC���6CQ��>������?�d�
�Y�?��׿I]�`hi���L�EM�}�=8�W�����<�����'ښ��5;cݫ����yq�V��t/��FD4�xu��
�.�&`FGul�B�G�R�� �����g�w$�9���¿\?��ڭk�3�w��;{�KCuXDBهe1@l���ť���ɕ�6d,��n��B񀂏|��*et���fAׂZqg>e�W��u�usf��J{+YT�Ĩj�������4�8���d��𐀃��	��u����M�����EF
�lk��<�y���`�6�D~M�W����U(0ƾ��R b�ߓ���x�c���j�rl�s����*�ch�{����g�:����.1N��������]J/
�r�,'�$��;�?J�%ӧ��n*�GA�������x�ƵM�ڲ�@����.t)^�f��y��{��y@́fE`��G#u��&��^m���s�Fr�Ś�58ϵ��s���D��ì�����t�����A�z]�׊U��n�~&����r����X�vB�KB����Rw�}�.���D*��3�?�l�u0�!!�l������DQ��k"�G�OB(������|6���g���i�Bc3�Q*\:Z�)#j�L�����ǅ?�j���#�\�����A�V:� ��Q�0���Z#����.�E�2���EO��ٺ�I����ۿ/�A_޿e�慳��}{Y����A����<�Wie�V�S��"4��Ḅ���?	|^�Ol��Q;/��n�t��a@%[1�>*������еq�������m-Ѐ��}˄`��ڝ˃ݰۓ:SV���Øs5�K�=��h%��j�[(�ǵ* h�T- P�1�hxaT]�+I}����Y�_h/l7l�-��;����w�R�`�I^dT'�@���i����F�D��X�:abr� =���׊a����q�l
��|��Ġ�A*��Db]�{��?뱝X/�d��a�ߐ���8V�n�j᫁�f�n߭^~��&�H"�� ���q� �
��dpXǏ��E�Z�@7w,lL�gV<z��Y����2�d�5`�o�À8њM>5��oƜ��i�'d:s]'��_QqJ\�g�A0�O��e{Km�q�7���VvI9yy���XB�mˇBB�x�#U���j�*�8;T �]�E���\�b�֧�6+sd˵�	�+y`BT�� Q���4�JiWu�$t�����Dڲ/^N�����:���dk;u�_I��@�P�������Zi7��:��ڋ�~�v/�p��^��k�8�̷�2�O/��h�ǭ��GFb�-�w�^�M#
��@+���K��h%k~����g5({�
���@ @�N�O�4���_2r�ܜnagx~�ٌI�P�E�"�̤̄V*���Rj�������.$���~ir���y���[�l:U��M�Q�%�~�*�BǹB��zݕ�|���X�4�8�ā�^��� ���m��v߅�[K̓��T�cI�1,X�1�Ee�6|�94�*aJ��9Y]*�*���?��pe׏�~�_ʈ̓�ՙ0#�3�,7�(7{?�D�3 ���nS1=#�zt��W/(���&�dw( �q�������Į{�<u4.������{�NCi?�V��yQ�vܔ��Kg[=('%��N z�pR�@ݝ��������>@ͳ/ ���~����I�	�;�V���B�=��гF���J_�m��4Y�F������r6�+e�Ę$�� �C#G�o����`�An�+�kL�Ŝ�� �37�� p�"��ޞ�󳚺A���8�=w�  �&�;�c�%����Hq�(�[V'|�\�7(�ޠAmi��h���)���"�@2.��С�P ��˚��,v�R2%�R�Ǵ4\�\+���8-�k�"�tKN�E|����9aձ��=s��Oa�; |gv-rÊ�Ds�!E%�D�o� �ߤ:K$��������s�q�Ň�Ӈ���v�IGB���0sY�ư�������cK��T�?�|I%M-�eLϔ�u�T�{�>��I�|u�S����TQ]	:UV{KS�-�\�Tl�E�8�fL�i��s���-��UL8�m]��m�g�? ��P���Z��'��O�՘}V���P��5�R��8�K��=����藋�Z�E����Wy�K#/2~����O�7��D�	��,���=�M7�����"�mu�X��ҷ��G�F�Q2�!��P2��"GO��p5���.>!s,���.%�o�� 9�ar/k�y���� ���fgn`�BX�E.��P��!^=�F��m�<�Ý���i��?@D������ �8��Jd�P(��N���V&��x�7�	���#��}Nl�����O�@�t%K�.gH�mŊ ��~��尮j�-�dd�t�]�&)��/GH��)yODֳ�y>5r�o�~K�ʉK]v�@̰��F�0���b�E�@y��N����jz�m[k�I�I<����.��n9����t�Rz���[�&$i��*�w��*岁HV��٠+E��o+iS�8�0Ԫ�� ��/��POF8�ڕ6���xƣo}��9��U���w�MC%.$�mO73B�0�Q&l�Z�"fD�B��j�ɸx�Mި�f!Փ�ў\Qވ�;3�H��.T���<6/�|�G>&�8�f��n,d�m�����5޾7�l.'�M�ù�礕sJ�NQ�s�jU}��"ul�Bt��穵��5��f�Sk�社�B�:nH�X;�`��� �6�\֕�L�탍N/�u�Ⱦ�k=�A!�Һ��~����eP ��6hCz�^����dVL�t��Ӹ���*TXF"e�!P���2+qp���i��R�+��X��� ���u�"Y�Q�Q�kkk�WO��?`9ψ����O�� ��\�ä����5Ȓ�]^�{�ao�ק,�vm^NzTkOE�ژJ�L�~�,6="�VD$���P���Cfg^��ۑ�,�[1���Ϻ�c�U��������Oh���׊�����/�ʢ�DB�������
V�H��S���w�3f��\�¯�m�L`/@�3^=��Û���U�r�[�o[3G���� ���◸4�E��ģ������B^�CnN�v�q�nyw�D�P2{�r �QS�"G�����<m��Ѭ}��*"� ���t���<��;P�X�S�%���+qz �[Uz�5��/���_��&�\O8��q��~�����T����2����ݵ*7��}d ��xE��C���oB^������Ֆ�H������=G����`�Y_�>5W��`�V
�}ap�?u�3��yQ�;�m8��| >���ܽl`������#H�<��Y�ۦW��~x�`�VF;��2�+�V�E�ZO��:��c^XX����|� �yZ���'��#���F�����"4􌠡��yfL�]��+]���4�I�d$ ��p@�*��S�H�\��~~�1�1��g����;m���	�$!�/ċo�X(o1`F����^�|k��h���&l�:�D΅�A�1�"G�.�.�H�שdN��y�����&+ka9��損�<:��w�k���։��&�����g6���y�kP�.l�hQ�2�M�-�Z�:��-�9�,� ��h�3I�k2r̯�/\���>�;�/�>Yy�I�Q��T�ݩ��B٩E�ݮE'��{u'ܮ�=
�^2C��=p�؅)���,�u]��j*�k��ʧ�R���=rP8���w�x� �&�3�=�|Ÿ44*�Dm�b�O����\��T��4�%�"���[	z�޵�Aϫ���V�d�'�&ewG��z�곤�}W7�	���@Jg'�pN|�J�{>H"��~Ř!W�W��:aU�
�*.��ץ��@��qDs;���H�<��_ 5L��Q9H:0	�O�+ԥ�KV�����\u�m�ST+��
�������W�M+�c5z� 0m���I�L����z��-���&�w�W��d��[-k�[���^�H�V]5z��Sf-\ea����X��2��6������!���ŭ=�[��\:	+�S(���y������ZB�Y^Tӵ|;}kE��Tp�-?��{(�N��ډٷd���`��������^�㈄��ݥ�z�O	T�߮���:�P�8����ZϞ������I��͋k�^�y>�C��W-\�t��:o[]�dr�C�.US��l����z��ɣB�x�?�f�Uy�5�m�RL��p���������Fd�+��~���L���?�+F�}�÷^�i0� 
Z�+���yͪ���X-��0�~���<��F�UP�l�̺��x�������kH�\��w��� xK�e�ǆ_V�]'���NC���w��+�u����tX��)�� �E��a����>�Q�����e:�a(G��A�|���ky��a���)���^%p;�D�R�B�6.b��>��@G�}�نܩ�4�M��N-�,�z$O�����'su��J���zY��sq�"����}D�]t�� �H���H��W�[�33e�fjp�{�x�Cmo�P���%�(J�#�*��2�	�+�E���Ho�ܭ�����a:Xv"f�+1�t�����!AC�ry�k��:1�ѽ�M�R�):�^}�3�46�\�n|@2D��0���kQb��b���gh�t��rL?�h��IC�����X��&���\ �fB����՝��|=:�aH�S�{&�L�GGL@0�ާM�ۢ������q���c�"���u\Fb��ci0�@b�iUs@<��4�%����a7��j��k�E��7%�����J[,s�;�M�Eh��]W����C �fK�0�Zg+��:3�כ,���Q=k	�>��nb�4/7�P���oHO��aE3���Oږ�k�T��]�{�:������f�`������1
��!�<Q���Pj�@*�IK%Ϻ�v����]ǀK�����k��W�;���^�C������B��
��ȁ;a_s~��\�oi��Z���;Ӽp���U�4P[����?N�3ei�O��R8z@�[<S��V�Q��4]A����� 		���u)����e�y�����ƞ	+|5y�I%[���^��u�?��TS�=*�S�������s]��|f�%��x�(��_"��o���;}뢽�����Z����F�nmG�xڹ�H�Ң�� O����RP������s{v��a�(!�����/�� G�,�5���r��ƌK��'x
��Dq�@�%̕����"�E.�7())���D��{�N�m�ӺX[�K '�;��/		k�L�p*8#FեSU��%�p��8�9^��햛��h��X'؄M@@�����G���/ON�f��I�PDOqZ�E�󉕽��>r����9s,��&o��|CK��M��M0}�Ж0�l2C a楑e�:$g����:�������a�N����A��� �x#-8��~U����h��m @/����k?�7�o���|���f�n��Ix �eF~�ŷp�Ϥ0;��\�K�?U����è'�-|�~��� �V�莯y�[Zښ}�%)N7խ����������+�[��6��D�0ǰ�ѹ��s�5V���C��
����~a%��2��LkT��O��{@Az+��~�����p��r�b�,�-��ŸF,�����l���H���'d�����c�����-�*�ݐk�n<��7�`C��U7���k�4�")>�[�BOJ�U��Ѿk��ÄAnB���F�ⶬ������Yc�Ȇa����� ��[Kd����h�DCR��2��L��ݱv-3�	[�y�G�\z� "��N��k[�j�_Ӷ<���Z�rE��L4~ȧ7�U} {���9�I5��9���.��C�;ػ�]%��~AFQ3�Ea?<gH����\�-�Gxo ��ރS� 
:]XT�����qo�`�1����'�w�wZ�
=�
��e�	�z�T߉"=�7  }=ɔ4LQ��,��چI��]�f%@�j��%�ߩr\�//�p'(�3��L1@(��Hi�`$�5�Ѐ��{eY'w���<��'v�NG5cFPpN�����VX�ϫD�����X��#�y�|���"�12Α <�kB��M����7x␨��p~K	R�7H�R�L�1��v#r�B�U���K^}+��G*C:T�t��baA4a#7^'!/W_�-sv�����h�j�3�%�Ƈ3�e�5+s�!�E��JS,�b�v��L�(�}��j�	�rݶȱ�5/�?���Z�U�t��O��☼��l�G��UZj� h�!z����4O8�#ݯ��]��h�<�"��+��-��cB-�tpX�R�f���~<�i�<*��`��&���69o���lh���}i�5S}���(�V���kc)y{U1�o�[���ט���˝,�5Sk�-��b�K����/���'�%�'��Z�=k=k��Lγ�Y���^HXsF� ��M�n�Rɸ�â�2L���+墭��Ph�ҿ�6����q��"	e��r�D]�h1E;��l�I;/�c7T�f`.�:*e�� ��������W��
]F�_In�����ݨW-Vv�_i������T��o�.W?���kٿ�y�a�2ԇ���J%W��o��7��V��Z{��c�G��@(�S����@s����� ��NE����b�v�ȳ�1Br�]F'o���8�+�p��p���:�IBvL�����(}Iq1��/��>�-*�% j��$�Waɒ��O������g����@H��( ��)z�&'��2���KI���v-�N�9�Ҿa�]�9��I��k�"t����]��R{�����uc��@8�|�4��v�����J%q��`��l����+�{��KKap �����P����SrцK�e2�7��4���wyF�]�/�W�+ƣ�?��u��jڟ��#)95���+����W1,z+ɏ���N����W�r��i���{�' ahwc��#�(vJ	n`Q7�"p��S�h���׻qnQ#����_,�lyhP%M0�ɮ��gB����U^u��ŃB����V;&��e�c����:�C
)��<W���gxs8����P���f�BD�%��в�y���mB��S[<Z���%��������;#�����蒙 ���t�Q�7�N�*�,f��͕y���`��C�c�N	�!��U���P��'Sc%�����	�ŐY!��(��Y����@��tv�r��j&���1��~�S*;��0W<��=u�P���g����˚�Q)卨����_�ݘ;�Z���~���!�"_Ά�_�4�n$5�����Ƈj����a��4}�{D/;�}*�8X��wO?�,7䠂Н��z��E%x�V�m��P�$������_`�o(���� ��L^���g�N�L}��Vj��b�b���8PBbaT3��L���6I�BYS�G�TS��F��ň�~����E2aTlo)#l%���v��X}OB�L��H�A*_��s�6�6��uO�S�2���"Ғ���lfhi���=���$�u[��혽%��B��v��Na��k���H϶����+�֨���jG�t�9\=�x���z,�W���6u?]����UI�)�p[�c��_(��C�c����S�L]��\�	T��r>���{a�"�ϒͫ��C�������,�z���-���9�$��%��!���wG��J�Z�����>���+�u���'��\q{[K�1տ� j'V-m����N��#Y�H���h)�����sm�B?�C�*�[���% Wak`��9T'�7U�M;i�����Z��E��2�t:��L�W*#�t+�y�xf���������|=[�1�����kF����q�~��$�ׇ�W�5c��P�;��ѻ�	oD>1�jt�M�aFc'v%9�V��-&��V������Yև�	����<Ge\f�bN�<VbL����Sk��P�N6�眬��Dk���E8m���*a��������2dQ�5�{�,z[���ʣ�}:o��x�R���O�;��2]�j����uu�n��#BN����O�d��}Lt����pG1�D�U<���}e�^�?/���
).xo�1;_"Mv`�c�����l��PW�^⺾���W�CZX��r��ʦ�3ц�b�]>	XV��j����6�Z�WB��{���<�T�5,�>���n����Q��0��s��|^�&��,�u!U2/:6W��D�/��a�|�a�L���D܋ŜV��T�j�U���g�y�\yn�5��"����L�u��� U�Q�%��Q��nLE���i4n�yG�(l��VoZ��=�ҳ�����g�$~Px���z{1M��$��x��u7�:vg=��ʝ'���<�O,��������%�|#�8�O���K*p��A���Gg�b����G��̾�A͞d-"�µ�屯���0��?�K	������@����׉��V��P�����5�$w|�W�=Il�O�lVm�XM��j�
t�U����d5����.\�G\���6IvL�p�uy��I�	�a�c�-xh43\D������"K�:1>�lY����Omn�̛y�M�i�g��ݞ�R��H���p<oT6L���B�켤�\ ~�f2�%�S�3�v��6��~"g$�bo���>����
I���g�Ӛ- �l����6h/���> �6�/�E�<�|�u�TO�aR*E�NԑtF�VZ$��)�gP��y���;{ı$��l�Di��[����{gT�-k>��")u��dm�`�-����2SwBRw�Kt��"NN�� xƩR�]����P�}n�~N%I|��\��{�^�ٞp�=�U_z�����rJb����G��A�r��I�XDHm&�^\�ƙ8ڶ���-�����/�������/�VÕ�u���^#����g����y1�4�:�=Җ�B{��Al~�	�4��=��S:7�܇�c4����$�\z��z�oeeh4^U�,r��)�%i�+�Σ��%Ԥu�4ᨫ+�	��, Z�2�<,�$lrD~������@v�,��V)?��V{��~6�_�u9=@7U�Q t�Dn���g�kz&}�-�	˭�������o��B+j�+�0�+�B�H:�ؤ���pRs3��B����2��ʁ?\	�SS#��\���٩�a�2	�bV�_(l�
���c��_����;���v���H*�x���12���X/l_z�=C����s7�S�}y� �fu��TVV��ml����8@��j�ܜ	a��%ob��n8���e6j҇���z�q�;Q�2����>6+(��ܑJJ[�G
F7E���<�@�����r�6D��up�9�+7Y��y� ��D�s����=
t�c��փ�)�F'����ǟ�+�wE��5�e,n��7����qe��s�.��ԗp�B��[�H�cQ}h��9P�fÒ�y����T�z�����\GD��n]|t�rH04�;|��s���F~m�n.dd������XB���"��LMM?yBB����+�ypd������ﭫ�Z}rՅ��#����h�W��n���n�:6�n6�7U��3l��L�3���{�q��Pp|����]�t1,G%��r�`~�J�)��ݬD[eN�e�]�JV9'����g��N�����R�� �/+nZq?�&�����AK��55�n��C����T�..ʷ_�m}��pp�:�=�٫��v� S]��#�1��d�E-4X�
H���i$���>����x��>���]i;��R������:D㠽�1b�p_�bo�3u��)��F�NYX�L3W�����D]�W��ƾmBu\�-;�xc��%���GI-I�ĠLW����������ͦ�s�����b^�����<F���:��m��TbXl�ar�eG�Ӟ)ܜ3䋋��y�b�����귃Ҷ����s�/�]N�֬."�e�����w�RJ�~�������.�b,�t��s��1s�bU��e D�at��(�NCL����=y���=���<��Ν����_T�^L4�������f��Pl�e�QC��� ���M��[v�E������~d��(�I��<=���m�g�;$���.��f=mu�R��̙��	o���N�|�� � *�OA3���7s������,���b�քȏg�[n�7{�����h�K�f�R��xh`�Ƣ͸���k���3m��������:�����ю�Hӑ�_�}Z�~���7W���o��粎��=|��#2ډ+ѧ�X���y.�]��*$|'jM�<`~twr�o̍���o�AQ�D�١���O���Q,z��m!��#�K�+��5&IP�#�����a{�6XR�󠟑Œ'��!HLZ�/WI�������s���uD��_�O�i�U3\Q,}���K1�R��W�??���;R�'���pך�Y|�Ia&ȁ�a�s�>+=U_����ˡ䀪���.�Ji>��f���<�0p�u��玒�R�~��!3��GR��[�%�N%�]��%����������H\=]����0���������`\����{�DN�B�H�`B=�+���X�w�q�:�&{&�)L�=�D#�����W4��x��B�j�?�͹f'��eV0��M�w�+)�/�9������"l�u
y|���xBC�Ňh�U�

�Al��ܐ����X��	#P����Ӷ/�����O� =�sz.f��FCP����c}4�Ivq\�f�ow?	_�v=>�I����$����T�X�%`.3��5��-Xq���Q�> ����1]~�h�@�i��9��y�8���zi֬�_�-��xL� ,/���$����B��G�>C�z
r��aK}��[A���O��µ�w�"*��I"���eO�B���k<�u����� �o4�9�H��o��4\ʎ|����7X@IGpc1Cܱٴ������5|���:��-�)+���SR���?�@#�z:�e0�S�^�%���q*��W
���l��fҐ7�8R�:/^&q��k����|��5��~f�a��%�3J������ń���jZ�8q2��!#b����Tg�SV��'�r���Ųԣ�c����8;��J�﬩o�J��Tt�noQͬ�/�~�󝋽�?OD[����bz�4��a�hYN$(��fQ
h��<��Ѡe�"��C�����#���������"�,�𱰘�`���ս�b�[��wuv�dv����d�p�m����6�R_���4u�Q_:J�9�ɀÙF�F˘:�'����^�5�
�xV��J�]Z+6��U�04�@y�:�T��O���*k �Ѝ�:@�`���c37�|�h}�pA�+���A<���m�3�t�o�������q�Xo�m�B;�u1�׭�0�X��뭶9koq�Z'UcԲ�K<���`r
�wNh�i�����5=9�G��r�z`j}g�A	����fv��t�/ '5z�KI=߱�2;�1��U;��R��x��r��9Y#����1̳�8$���z��8��b��秏�܀�����ʷ��E��<�w����dti��@e��U���7꧚�1�p�����*L�-���*^�<��ks ~�\���[��c���HG� �1J`��oo�"c���۶�h��G�W����Ws���;�)!��x?���,M��Y��Vl��KU�aw��g��7�Z6�Q8������m��̶����@�����f��,�:��l�S�]�{�W���~|�~$'%�]�+Ќ!��t�0���l�����8��F�Țo�w���(�#_N���~���Ǘ?�`H�徜����66���,�,�'��ܮr�}Z���ї�ॎw�<�ߖ���/V����hD�3��[lkk�g�C��~>����(�Z�~	o��cV���������l%�\Q�5x�?��Ϗ*��
_���I�����bN���Q��2~�#
㰷���(1��������è9�U��wiY��?�ҧ��qa��h�))���;���jC?��z�'��F��?��Qzyz0}��������9�#L�לR��5t���x�� �_�Y�G�i���)�i#[���}
�L�uGM���ٰ4c��J�u*�O�tT��ym�)����Tj|��������
�и�x�7 T���S��V�ШԲI?�+��W"��{��_��s�X�G�U�K�gwj=�\Z���m��(c���!N5�t>d��R���j�p�6JN�y�¹�1�f��'�^�$_sSE��p�r�S!�(M����>���D���"\���Gc��>L}8;�������r��D���.y'�F�־Ƨ�!�����G�`�;��S*��q��#F��H�8�`��e�v(�����(`���Mғ�x�:�B	��#�E(����	p��L��JL�����'�VGIr]�8�ќ�hr�C�3��6��(�[y�����'�������mr�������ZU��˧z�h"Wvؘ�T��()ȏ���d�"�@;㿳W����e)�;��D��"��1��|�~a�����Y�^����?���4�n�q���N�+�a�!I�(c\^�FrF��GdN�=��O-=F����P��rb���4㷬O�|��C���Cc,I��- �ڴ�S�>���d:�~���t���[�E�}��<*�" ��4�"݊���� Jw�*"�H7H�  1� 0tw�=8��������z���k.Μ��^{��}��7����B������~�>��İ���@��&��Ap駏h�o�턄$5�z��q~�/�'������-,q�Q��6������?��.���o�!�1,X��^ ���'�[ހ���������C��=�$<p�����I�7J��]5}%1L�����K㽋E&My��^|Ry�2��j�zA���%�މ�5d]oZ`�?ْ4�ш�J�oc8�^��������������y��8q�g��5���6'�G�a F�W,ĵ�����3LX9��7�*so������HH�묄�.�UМ�5"�����QL�x/c8��辊#��]RU�U�h�>�����s��DF��� ���ܴ�I+IX|��I�ss��c�G���#׎�)��������@^e7��]��}��"�g-[�i�՛�(�*䆧�ʝ(S��Ii��~>�ͤ -�����7�*��k����ױ��%�̵�DD��l��yd�2���ԙ�]�/�ڿ���󳋄�G�+��]2;��9a"�ϤZZB�A�$��TR=�RuBfao�+���$H ��<�6q�I��&ٶ?-+I�cfF����$�G.*Bu�۬�h��dibM����1�Z&���h�ϝ�ů%{Ẑ���٤�C��s��J�X��ĕ����Y �rG��-}K��0 ���׎�5��[b�������X~��;���p-�2tMp',�J{�+=�w��z"/����hh�e��s��r)�:D��;���Ƨ˒9�D5B���B�#nE�)ǽ�E8m��\�����k:Op��,T
?ᬒ0��S�8��mi�-y&�p���1%�$�l���3FUm.r� �|����|�=N��i�G�`a����z�ڷ��S�H_
�;3�4�RH��E�K��t�ʌ���mu�{<�#�G�Xx�˼-#�R�����۫��9g��N?9�����r�mMgcz��,b0dvT�Ǖ-�M��d$����刬V�y56 �0��X"���x3����VW���v4"�#+:���ܥ�I�w�R}Ga�:J i�jE��;���	yl,U�3`�:pU���D����r�%3 ��n޼i�����M1XMnB�U�,��ő���F���C�_;I:��1�$���v?>�7�Q2`��3�m;x��`B�ĩ��1�=N#a�;'�@{�ˈ����&	�JX��@��$[ae��9Z�������
��WY�
�Sm!]+pR�d�6f��|���#֧�+.0�xEu6��y�����*9��W~�F�F�K�\��q����(˔J��EU���5���BF�Y�Tо�Q�Yr2����ty�O-��~ �h����M	9<�8vjCC�\���k��B�J��0�JYcccWyGGG���������v����Gz�R����T�k�h�jq{����S�M;��z�z?��-���L�&��8N���6G�#z,�?����
?B�p�����߾}�{����e>0��f���"ҟ&B���U^^��DFQ��3	{]\�*c����u��1**!�^���d��d9ee<���>���ZaCM�����?�\����?��:�����_����]=Q�����A��[�����Y �;�hy��bG�q�[Q�H��q'���t9�1��"����N-��?<}�Z�Z�Aub�L��;F����|)�sx�\�J<��d���.���L������W�w<XX#C�m��($��#1Y�������Ѵ�N�����J�lz�]/�T��-f�F�w�������h�n�JM��r����D�<t
���k
���K������
�݌���Bf��uT���F�;]?kn�i���{0p)��F�m��*$����/���3"t��p=�tx�4&���ᖯ�s !Ӓ�H't��|6���*�T0)&��
(v�.�Ѿ���ȡ�@�t,�LOttP���>ǻ��⣝"�h�D��_��(��-or�m��f����Q�=q������D�h��Ҍ�j��0�r�=V�<��I�MG��jT��2�dB؈��Cf��b?�K~�*�lT�yML�1� �����5�;ۢ_��A�K��iC�����3�r�그��9R�m�dqt�u�;��h	 �X�Xz^FO�x�c�p���\nٞ���v�[8��`���4���G��Բ#�����g�m�}�����`l�Bč?*#
HM��rPSk�BG�������a\5M�Wyu�^�g~��T/��t[�ød�P��e�^d�_CqM�uz?C®?����^����}񹬛�펗&1m���ۧƒ�)ĻM����	/��[[l��~v�NT��T%��G1�#/i�ao6�f�m�^G��<�LV�Z��;<�b	ȋ��]V�Lړ�T�:�'�L�Bf���A�գ�6�y?�̮�f�:�wT
���L+b�to��'�4�7�|�-����p厳��W/���~f�Z@�񎳏�<xi�g�;���0�Χ����h{
)��8+�wI����"P���gGm��-�Kc����u�ழ��!��H�E��e���v���

�kQs��k1L�����1]{G�ſ���I�g��5��o}����f:V�����5�&�$����h&B��G<���.�V�R.���U��˒#f������3���ۤ�v6 /��z�TM�}gD�"�����s�}�|uz���o�?�ž��S�K�@�Y�H��v�|�τq��R�gE��B�'�:����'Бը��_���tJ¥.Q��)�\kC!���]Qm_����6���O틀����V��\��8:S�贫�_X���4�	K�7�gkur���w�-�a�Ӈk����p�T2�aS�P���֯�J�Di:B�"�%�:e "1|�pH����3.Z��fT�11�{M�t��őq�Da6���"���ؤ�{������ԧ����!�i1p������;ܨ�zo����r�������������C��
> �a|�azU���N�>g��-Q���f��|6 �z�Hz�]y�(id�h��U���Gs{2���S���Ŀ~(��_���l���rb6M��աe�s"}�G����=�
'���R[�,�fV���)U�/f�&���hlH�n�`������!�B�T%�wdba�
]Un �����ll�
ϝ����xH��ȭ��"�7r	>��s��d�/��<f�qY4&�#�,]���|2���G��\i�3�A&�9?����7����!��]���5�C�h\����~aAK��X��>�� ������TS��g2"����e�~	*��~_\���^��a�H�\���"�KX��D��3�L4Kvx[XJ(jR�ꓞ% �4
���մ�X�}�V����q�A!7#��h�
�Iޯ1m$��&��{#g��yt�\2-�Y�R�dvo�ų���8���GE{���Aݑ|M��� |�?�z\xm�|-�g#}�	��#Ñ���_�p�k/0�Ӳ9ټ}XO*
�v�I��&��W��B�rY�f}QW�IO�c�ֲ$Z����Jͤy�����pp������S�|�l�P���A��@����-�/z��*M*;�l�����ဗ�\�MCT�^`���v;����DG���T��t�t�41!��6����y�-g�,��<�y��s��+�^

���𹹨�j�������C%�Ʉ/�}�.�ב��q'�7.[���$�#�Z����l�/Γ�O�8��[� b��K�̳���<CTy~���^%�f��)^%T���cȫQSGF&���"��T���ո�=���ہ�!�����ϔI�M��L�k����&[|e��~0�_n;؅rI{��]S,��v�|f|�a�[[����sq�װJ[����"����ˌNf�~?5 ���GJ>=����{�-T�
�����cO%���5��c}�����5(󷯡�� ��	;L!Ǫu�?7��}�FeζC.^a&qk�������R�<[���PE_���8�O��t�-���C�v�3�8:����\.ڗ���.�{�UyS^�(�cN_Q���\��ݴ>�[�侄C�s@��M�+��I%����&�222���@�v}��o9�` +��مL@a�[�܏�
;��Q�%�7y������Sh	<$$D�x�5�b���;����v%�#�
�+h�0"F�Ge�3寈�Cphi����{:E�z�#Dg�o�ť{��t^���É�x4!!j;<x�"`�� �z<k���_=�2>?2�l��q�����ņ���@�Ʋ;�����^+J�+�/4R���%���)��5΍�q� {F�=�"�7��_G�.��ݓ@Ux��jQ��>�-D'N�{y�ڎ��i4[ L�8�L|��-�7�T�ik�sk�v)c%�A!����g`�o�=���Ѩ���_/�:�	8?9^\��p�8�وZnz���9k�������~¨+��`�0!�y��x�&-��-zĴ��X�N��}�D>]���{u��h9F�4Kށ�~-9k�_��@���6�sm�(�`d@V�uJ"��I���㷸:Gt��n�wDH��iP��ױ��#��\���zz��V����%���X�J2�r�=._[�n�/.�"�p���ˍ�h��B�btd���	j������ꇳTV�
�@��QI
��Z���	�;���#(¡���,EU��� �g=��<і���{��Q�֒��C��K�|�H���|��Z��{,U�xNa8�Qgܿt<Awes����Y��\4�B���e�h��M���)ů��� �G�n��y5���9�]����ҏ=�R����{��!��Ѝ���1	攺l���b����K���ѦZ/�YTq �:ef�X�I箫��l��XU���|�9�P���W�H��N��5�jZP�y���B�z���mw��n}�t�*u����r��ј��O��Q��*�4�O5�}���P��b_��#�����u<�Ŭ-I���fwk�y>6.�ڧ���z\��JW��$Դ's>d��hI�������NN�m���V�7�8�=�3�_��a���'qDԲ#�gR<䭨���^�:D��S���ٟ0�xƄalMf����XT��{ۚ�N���v�� r}��gmQ�K�� H�߱h��j�A�:�ä�ƮqA�/�v���� �9��l�� �Z%68�*��+}X����J�P��5�M��M��#3K���bS�G��������9dGj���d@�Y��[wF��;��%�jV;p�vD]�7F�C���6���l��'�i��ю��v�f$)j|f\.&��+Si��9�vK�B=ζj����t"�}@�ۅ�O+j :���h �1����������.Ω	�\�y��j����z�!u�Q|�l�̙��!y<ƚz�oM��tܥ�����wz��N�x��������vL����U�1�fk�&���D��G����)J�J��:�RZ*�)�������iPe��Z�50��� �����b�o^��aX�<tn�^��Dxu�� 9m���X.��xuO����܆���q]���	����+S�c@��q'�A��ʿ�y�ݸ����a�3!�m��Yj�Rx��3���Z�f ��_Mǎ�� F����Ym�a�m ��A5#t!�rq�\��ּ�c���"�����\ ����,���K譄vGc*)���u���� _�T���ZXRR������."2<��aʏ<����-����f�t���ϔ�6�iPe��c�e��?��=�7-�PЯ���ʥ�����_0{���}_�#m%�B�C�s����㖙��[&O�Ofb�����o'%�WNW�
��HT��c���M����=aaoѥ.��t���UR�/{7�u�~��g�~��k4,�
�x���`�vdNN�Ygh��5�/R՜v��__n��y�U�j����h�j[B�r��.��x�z���/��iUY^x��ã]�v�~���kTg �\����W�=iX{��i:��<>���oO�]���S��gz�6f u�D|������3���?i��}v��������S��z ���
ћP��͠��ɚLD��0��s��T�'�䴥
A#Z�2���ٌ�U������\&c�i�Wiy���g���L�+\eWgtW9�p�"�a���;)��#�r �ED���S.w�u�a�+i$�+QckG��n{�2CN �8���G �2C�(����^�&v ������3����2���D>�z N�%	3�7j�0Ѽ�4_i���Sq�]ݨYM�g�AO7_���aa�x)��sz��3q����DF�*R�$����woc�\i�߭0��FI̖�p�G[�ƩsN��\�:��=���k&��ɞ��Y�ᎎ��U䖪�X�z����e^�/�N���b$?o�����]���mm��<(3 ��ֻ8c�b�N�Nxه�d�V��A�n�/U ��XH^���`�̯��ltep<��� �9,IpV��u��Xu+#��D�z?;��3�!��w�B&=��b�l�Az�J�{�G+Ŗ��.��FUv�}�� m *!$������K��W��3��Y�Fbˮ4�r���c�%�/���Q��Lmp^�x���l�ۧcZ���L;�ve��s�bc!$F��?+�m�(T��u	����`��'6wI9��e=����ջ�rb�?��&���H�[�0�|q�U�jKO�2�c� ��1Jǖר0�*�el�@;����K��l&mb�	ϒf^%)�/�X(��� I�X[swl��
ֲ�X�k�I��������0{�ظ�٨��Ŧ�]v3.��:F@q['l�
�Ť&�Aa�_+�R��]y��D�R�f���@4b�&2dD��e�a[f\t�cP�=����^4Q����鄛h@��S�+�������D��'ek&��#���?g�׾C���H8x?�e�4���@�$`�E�D+��zO ���
Wߟ\�S�߸��Z&�0Q&ĥ�@��W}��6a��O.��NQ�.;e���j}w�pc?��^�b^O���C�C}�By�P���F|uɣ�Ȝ*�:a�yHr,>�BTJ�Z(�3�!��d���7��d&t4VX��é����B��`�EM�ܾ{�[��3�a�hś�E�O��� ��G��Yi�w�׻�/�ڠ`H)�)2<�7�t��?p�N�I���K��y�c�/g�%ih�S�;�N�MQŎ�W��B���N}X�`:b�nȵ��zj��r�a�7��<���^�O�Is�����~6}�3OY�u���l[��������$�g䣌O��q��w�'����0�l�9��5�g�mCFxΘ45�,'f���Oq�p��-�\�!����{�d�˓`��X"����ca���_���0�Z���g����??Q�|Ջ|hxhkt*W��p�����4`�}�J8�:N��>�<--�妁J]�Z ��䈄� ��k�	q�V e���Č�N��c&���4K�� �IU�'<eX���PxK�퉂��I���x��B3&����Q?~n�F�'&h�|#tl'\��җ����@�Sb\܅n6q�׊uv�M|u���1�?J�U��Pr���H����{N�F%���(Ĥ���)7��N�JW�"�[�;)�|�B|b�뉤�8�����<*2Ĩ�|��O^5gZ^k+���з[u�\�)0ؘ��+<
�^Ё+��u��)sr���eQ?kwqU�����ay(lǴe�;��o��˥e�v�[ц�\C��m�А��ʀ���&p�m��sЫ��E�,��t?	cNx��2�ۻA;$ZQ��ȵ=
��Je�Yz1iӠsZ?������5���Ûu;�h�ff�ޏ� ճx��=U��Sp�g��떰G��.��M��٬Ra����hqyX�z�EVC̒�(����c!#�)��;�Yfq�Z��ǳ���@��j��^4pg'��L�M'<9ٴL�˩�īY���s)�d��2�v����gE���_�c�uko���4��Ia�x �də2GGHc
v0�pާ�b�S�i�m`C!@�f9�?$���=�lװ�ۍl$�ㅕN�s+,"I��<��9��w��?T��B\up��v=��M�{�'L�6�K�@k�q����j^0.����@a�������Qʲ�l�byހ��D�Poxf�z��I02T'��j ���}<Ã��GzW���jj����Ƙ>��}�q��Gl��Vn�)�]�v#�|���kA�٭��b7�,����̋k�������ʻ���Q*0�4e�J:����Y�{��g�W^Xq�@F5F���,E���ջo.�4���R���y8H�>L�=4��`��P�ơ?)�����=�$l��	Ku��B�΀�v���T�ӄZ�{U�-<R�<t�>��ܯW;�8TR��5(�z]S��>y�Ų��!�6.�6~C�~��w9��o]dg��,Vir��
(�E�t�P�*��/�|���]����@�p����T�f�N��w�qD%�oM=��n٧��y��f��OHj�X@t�J�e�܋�Y�����/�Y'�Gdŧ�n��7p�z=�8��@3[6�{ox�z�\mmEL��oA�Ï����b�B-αw�~㷻�J+�	{�*5ҡ�v��nёFJ� �E+$4H����&>�ڕA����sf��'n.�����K��&N��P��
s5yO��77�3ĉ�����8�,�hy��M	�@fu֞����r�;D'E�҃v��]�nT�0jۚJ�4ʶ��m4�Y�M�g}�ֹ�8�(�G ��L��O�J�7��g�S>�Ȧ��W䡙��-��b���Ct��e4������xu�e
��i�k���g�i}'��8#Rv4SF�؟]��^Z�����y[�U�{�`��@�_�������@����g�X�[�|#3��	VR�߾d��3=�x>�ڮ�Q�>�=�m~��0�(���S������blΦ)�6.ݑ�?�A���`ݱ����� �=p:uLC���sZ�N�5���s?a�v⸫�R͇Cl<�
�@A���7�����
n����V��.L3�udJz�74��v���_���O�
�c�{vFp���WdQ�;.'���	��z����\��DAr=k��U��>K�,�L�G�ȭ|����FJ 5n�7�$x��ΰ�QEM��������$yn��x�bg�&�K~��GOf�g��6H1�A>��k�-��䃶sή
���$�����D&^�"�G��L��Y�e:�
�q �ޛ��qC՟��2D;]҃]�!n�G>�&��V{dN)�HPbKPX��Ypx�i1��E��cN�R_�W>���N����wO�6��p����q������tj� ';�g�0���#���])�[�|o���Q2�`��/��=���6Hk�A����[��?L�Zdu�
���kI��*���������>\\g�O㏽�$�c�&0����0%�3F9=�M��q�'O˒M��m?O��79���X$���ri	1��nօ���p�wb�I�Ʀ��9NU$��)�H �,��鵢Ƣ��'�yRY�����S��q�f�֛��xX�e"/����˂s���w�=.�/O:з��_i���;�ұ�`�K�`t�)�*)�*�Y`!��Lof��_�_a�G�X
�r)��٠%UEM|A�zn��[2�i?�����Gs�
xTLB��L=�R�UH�t||`�,J��J�P���R��i�W=�~�3!/����Q�Zo.Qv��P��]GF��g^g>�@-3�ݪ�aR:$k�� ���@L�ވdY�0}Q(v�8��Ѩ/'U�nH���߂o����[�a!�Z��l2��8e�qØ���b,�+�T�!�Ds8�U�b����`%�_T��,�wS ?��Pf��V�V��l��y��G��x����B�(Y٨Se��[���,�K�
�3�ݸ'[��\ӓ�xR>/���|���K����a��7�����@,� �m�SL�8ڥМq݈O��h�е�U�H]������9�5�[��S�ۓ]&�s޹-�f( �\��"i��M_��Y���]��.Us�{gR�.V*�t����3�ۚμ�(���HDμP����-�x֬W�;��P@��,�ϫ!���e8m>g�xZM#�U}����f�'R�S��P����웓��N��~Fv�Jzz��?�a�z �!)��s�#Oq��:��Q������b��S�O��aT�@�����_��Y>c5�U���'>z��$ը��5p�/��"�x��ѷ/ɬ�4֐i��c��&�Ń�'��k|�,[y7��d��&^�wAϿp�0��䑵���x��Á�(�*
�ơ��<�g��0,-+?�̾&��)�=#�E���,�����lm,.>�iѬ�6���9D�V�t��Z���WX�|/���r%>�oL��o�JF�Y�	����	���P��io�m�>	N�,�(��~ ��uC|�}`	�%�,L��3���4%�"Ի���w�<De�v�t;�W�E����IRmTVO�?e^�P��,RF ��sY�G��dI>g%mi�vr�ħ;�N��E1\���L��TvM+T+��(@.[ؒ�����?�5]���.�V履��%a� _L�`��#g�D�x��Z�ޤ�z[^�7`t�+�Q�%��jU.f���O�~Wl�7�N��	�M?�AxL	o��F<�̕�0��X��wߝ��8���g:m�jr��}��[f�r�im���~>��%� �h�8U: ��_�G������M5d&�6_7	*�&�e�	����@f��}8�����s�:-hˑ#���.[��8*��ܷ�I���@��4����o�����I:M��/�1���)�k�%�6Ok(�RK;�}���/��$s�����NP,)�v���G>�բC���
g�v�v~���o�dHMM�C��U�<���^1�9٧�W&d�������	�]�}^�?DR2u����2�%�KPl��;R�=������e2B6{� �igv���5� B�Th�7�x�D$���ϗ��:�AF)R_/�8r���f����H�? Y�R�(᫳�㥵�W3%
�~�o}Q�w��|Wr�E����A���hX��y	�(�c��4j��0���ї���e���GV���dN.2�����2`�K�$��q�Z�¹V>�&�l�{�?�o�g�����G���76�h��y��W�㚭.yGE�OU^�9�(��"y�p�n��zL$ј���X[�B��?0x!������������ї�)sW��R�'�x�ǃ�Ky?'sLߞ���A�lR�X��e�~�d�����r���=/YX����ۥy�`���r`�~����v��O�YTL�a-}n	����(��� �Ƿ�+4����k
�I����qlǑr����$��rƿ�d��똄f�s*��Ч��D���@s�n��-<�r ���
���;cN-?�� 8D?����s�.�V�U�'���=	W�`� �vj�3n*֑���/?F�i�U:��Wg�g&����h�}��Iլq��~RR�Շ��U���b!5���'ձQ[]i���;D����Ja}��_��is�G=\}�B���ހs�]�MM�D�t���pJ�ds�k�o�$�G�nʏ�n��<o,�+H�������P�my�w�tV@Y�G'�'�wz�Of��{�F���ӕ⁠���[�tʯ|�'/`��#;��f|�5F�:��ac����������D��D����	N�c~~�xB�V��j}J�s@J��5T�����7�p�����+!��$��q#lkҚ[exl��X��ëR{"_��s�*q
lo�+��~X���z<�W�J0�Yc��f�F����?ֶ�/˅���.������.p�����[����n�U��.�A@0�6rV|2�q�ܿ@��׏���^�.D%`a��#�?�q����ɢ���G�����p�l߳��£Eb\7#�J���[s��׍|Z�dpzkpޏ_��
�s���M��A�/?�
B�=�Y�v\�[)�n	M���fc7%�b�'�0q»�x�R��S���E�A+]s^���Z��ߊ��t����������u�r3Qiy7ou�Ut�t)�џ1`�KYH��#�f�j1ﰛuI
�?Nu�Hr�TX�,�VQW`��|!��#�Z��N��vǤ�ר�×�
~��R�1az���/������������3�Q˴��9!�&�ǴX�N�娒���,N
	ցQ��&��3���O��8�2{ML����r0c�Y����M�Y}�3�.�Jrpݫ�`u���sz�U��(J�y�Վ0Q�:
��zu�~���Ͳ&,[<n�
����n��o� �K���5������%8�#xW�Tʤ:S�,��0э�BO��<&E;U�>�ֽ���Gb�f��oga����x�<B�%4���x��.�߹V+�����&�l�"e�NJn[����j���Y�-��a��y�Y�}83>��yr�����C���>r��Bt��s�Ĝ\Z��O������������9�EmG|�NO����[�L���є�z�����z��x�`Yױ}I�mr�\�Di�X���n��)�?=�B|�jL�pL��H��Ts�<�ciP�雳	��˪p�q���Ae<2ЩoE��_s���ν���\]v�I�V/ωi�0���[ӏ=�c��MJ-�+�e�Z 1+��V
������{�����	�Y�~�aQ�Y��R���CٔѨ�&>�����1x@_��]C�Y�2��Uۇj+B���l$0o 8<�]?���}W�}���C�:�`���Ic�_�u]ӕlC������Y��Fϡ0B���@PV���b����?���k��)J�^�)����'m&!�]T��E5A�R��Oz��3'�Q��՝n��ԡ�Y�,����Y��b�Ür�V�%��J~����d]M����"CfR)�5�w��R'��w;\�0P�c��Yxnu��N�=�.��i�W>����� l���P�
RFiG8���	*L5�Ҥ�8���O����'	I����ϓ�Y7O;�=&���HpH�h��r��;��ާ��m��b{��4��F�C�>>�1�Z?/l�F�����Yϧ����M��$)�+��y|��[��;��
w�9�fUA����^���B���+%���:��*��̲]��qc��9vy��'�߼z�5�9�W��ӽ@6�q�yT���� sw��\Vf�de��"H�������T��"���!v�U[�2(Ė�=0j%H�q�Fx�EY�^�B�e��:<a�R��@N\h�`"NΗ��fmUS�J�ۭ*^?�V/�+�$QĻt'H��������'�b�N��?��$�=!]NQ����l�x�<��ә��Q�
��m�w+�O 7L�3�A��gvĻ�S��fRT�ҕ�ٙ;L��&��J�Ȏ����YZ9Zj�2��L2��A�[:�H�����=2ر/���c-DBhD���q��}��|	s/r�!v�Z�X��G�����X�B�Hx���9�:�e:J��:���Q%���$�<�k|�v$,;DβŪ�IqM�Z���1����6\��)B�"�B�_;����C_�.2�Ŀk�;���p:_���w�xn��;;
���Me�wכT��dA�A�����
����?���?<�:�Pċ�S_MQ���jk����}
'~�L/� >|ӱ�/��6Q��G��R^gЛ�UD(��`��l���'h��0���QSҽ�c�<��5�1��acq�$����&���6�t���,��A���QQERŠ;������cd�_3d�M�z;07`�z-�}eɟq��r)���*e�&W�H��&���O�|x=&���P-G��l��9��0��,,IGnKVKV`�2z6�&����EQ�[N:���&���&�>��MDDe�E��?�C`��!0�!�G�K�i��:P�*��*dM5�[��[��	L�8lM8~J	R�rR�*����o6�3�:��y/}�&ڪ�'�?'|�f_�W%5������i�/�LR�}�;��M����'��wO��9�����������H ��\� T���I��b4�ߞ^����.�٨��i�L��"D�g0�y�-d�=��f���n휩�$\�^�n�O��[�`ٜ�Oڟt��X���f�y�A�=���Q���}�eV�eL��KWp�'��[ǻ�~W;ΆK1�2^1\�tc�EI�)��3�sIr#!r?���+ _��&�Iw�p�G2q(�+�O���@�801����x�$&[&�ސ�Ճ������߄�u��.��Ev|����G��=�J�o���X�@Q#�Q:K��k���U_���%u�t�t!�mF���C�$�T��n_#�a��}���,��~��e�����hO�پl|�H��-�[���-\,{��ⴶ��!8�ʸ���%����7��X���Y�킛{ }��{��:��Ց�'V[���6R,@#�7��������9�O�k�Or)�CK���X[��p}�ͮ�c}�̖U�y�����2�wE�V���=�e�a�ros��n�3`�u��*���)�j�t����#��JZ1 0IXӕ!���5<e?��MYp�^vӗ��VGT\<��M��g���}
����L�`�Q)��#���;//������y*&J�l�h�:�ΠZA"��hu-}M ?]�'ue�~���#*Q�REl�Ԥ>;�~/ƫ�g�Sr�+�m����d��
�,}��6�t*KUx��Ŏ�N��6=�py��|�Rc�g�W$�����p�u�
�(��S}ݺ�����D��
�z�ɠa�m����Ͼ2ٞ��\��M�6{�MHJ�]�ڼ��*���R]���S�X���˯+�r�)�A|6U�!)�R:��>b�u$���ٴv�����vܠw>��^ :V��k*(g_m�m�{n�r�ot�`߫�����[R,<�Ѕ!�b]!Ƕ�~w1m����֒ᐫe�	4?m3��k<B���Wy\��hO��R�F��z���;�U��RD���H�i�u���[�m��Lfŧ����|�֖�Jc�s����Cm��5�D݄��d�,��d��6�;/��d�}�b��g��.�====��ްS���i�(��<�6�+=tg��o����Ծ��k�mJ�5��6aSb6v(��E�ލ�e�Ci��UNž��`8H1ץ�����?�g��0skOz�C��蟃L�Հys�����ڟ��4�}��y�Wj��V8b�e�P%U��yM�-���I=K߆���HД�o�AJ��a������v�u�����n���u;S��/OR=��+�~��i3�j���᣿u1��P0��������aZ8��o8�U6�=L�~��7��R0?t�gg�Հ�rnY-�5˼�+���I�4@NFŅy�(U�-.��$��D��d�@��:�6�=�FY��c��M�Z��u@�>3��i�?>�wА96���i���0Xw�K���?>4�$B:[YATOx�IrC�%Iyav�U�=#M�J��e���b<d���ڇ�2��}p�njBph���:b��S'1��Mqyy%�t�ۡZ�qT\sq�~�0�B���Ɋ�8��T������v�y��7}�pwX�1�r�NP&P I�NT����gų�(SJ�ۘ"�宽���`�<���ޟ:b�5Ơ*�|�3����4�v�o�-	�v�Ձ���%�3��@�uՊi5髊�l!�����/�{IoY��=���H�5���Yr��b�OG���]GW9��Vܧ�xS*�L��nj�d/JY{�
�������G������\=Y�<?�19����Q���盂��J�>�8��D�םX7o*m�,l%Y���hl����B�L�V��f�d��ؗW�f��]6|~𼄯�m�ث�2>x0f�vY��:j���$t�E���Շ��{���M��{G������U��)�7��o�b��m)5�3�)��#{���3����И{���yS[^I���R$�m��5�
YY��x�J�Y�ՠ痐�?1��H�=㒃����?[��IG
�`�
T
����R�p�e��R2Q��Sց�LlPn��މ
��o�K*�iV�1-���Ǩ�����(��hG�B\S�B�%����^�E�#D�>>�[y��9w�˲Ԑ��7�Cise��U������O��&�k�V�rJi�-5�?���V�Y��ϤP�b���!�S�3j^�D�g�0�0�<'�*���q%5�\q�:����[k`3;Ŗ���YJc��2'n7(���˳hȨ���Ŗ��x��J�$`�S��� mކ����OL?�1?3Y�Ǧmv��nz��K* C�j&���s��Ҽg�q��L�}��P��h��Ns?�6i��7ߔ����5[���W}.�Hŉ&a�+Q�0Z���H�~bd����A����A%oY��L��R����4r�����=^t�P���a*[���e�����xE.=��٪6�Q���(ďF�˜�<��?��}�R>�~�L�-Stq ��	r�s_�h$]�]L!��w-�YO��,��#O��)]�������,������-��~��8ɕR��E��j���ȴkʾ%dp
q����������Y���i y��;v(�K�XVXW��$�J�L{cX���vM�j��ɶ'��dN:ٶ1�I��ɶm�5u���������u_{��֍��S�Ҍ�ԯ,�>�{тrd㰭�f���HM�� !ޯ���\Sl��ߖk=j��VY�\�^-+��l��%MI�z2���t˻�ee�G�I�4q��q3�ڢ�Z�m��DLk���o/?����O������z� 6G.ʕwW0�ޢ����?O_a��FY�%��~RZ�����m����%2���ӄ�~�8 9�_-��i]~p����Jgeť�����b�,�	)EY
8�<ml7^�`�h�s����_Ϲ�x>N��?5�����s<�yP9M�e�#���bsr�?�z�l
�t&�sns�/�!��<�9)�K��
�?�.k�AES���톫H�^�#�� ��_�Z��`��'�5��:�t47T����n�(�8*�i�[�r't�$��?�g+r7x��;�qWeYm�&i�qr�K^5;����o}�U_�	~�(Է$b2�����_,8Dj��Q-)3��Q4���[H�+��ɴ�s�,g
���g=� ��3{V�/����`�I۴��@f��z�E�^eN�P$�g!��Gѯ1�U���C�� !\̥1g�7��6����<hTJ��3��
dO8K�m�ռ}_�nˎ��������A�OdF��*0�q��p��I��Wz8?�pc����s�d�4�9`3l~�����-�?��mx$y0?�(#���j���t?�(�o���.gWe��:�u`(��벉8�:0��Z������������j��̔O���$	�����h�2;P��m���2Ź�*��)	�^��"*��	)�I�&F��3c5Й��b �7	֯�^:8�4ȍ���xB��|N��ȏ_g�u�c�u.a<@x������Qr�u����_{S�ͪ�O��v^�M�{穈��~=!��'|�-���<��8�㠳3��߅(�ɹ��tZR�٢$qkzB�m��M��{w��������"���K�s<^�	v���I�X�_�0�^���N�:�ς�Gv������N����ݫυs�N�u�?=ȥ�w���v�$e��8~�O*L���ND�nןc���A�CU��������)!7<Z!^@�[1c5m�P���Z���W�&'�;%�۴�g��� ����x�Q�o�2x_���'�����%�F���������ր	�DL�s�Y�,A�ߧ���Y%��S��T|ي?/=�M�ܲ���c�gt�6J7\�r�˾>�Y��J�AhM2�-(��L��Y��)<BQ]��|�x���[��a	��q7w��ȳäQ=at�c�$���FB�yL�)t���]��?�9�����^����f���M����m�Of�@�D�n�Z]��#����f�8A�w��~j�؁�I��=��}�>�cų8��﹔�.Z�����o#��ΐ���<�H�Z0��u��&{��";�}��f"��Bo���K�,Hd�ħ��Wr~�WlwB����&J�uϺ��%�|Z��)�t�j8�YQR�y�J"v(�C���]�ݗ	J��������S!�Ru��i�!�D��F���u	�p�蝬K�?��o����a?�����H \�y��������mWG��V4y.��Y�(en]�U����L��g��l��2��8����)T"�8���쵻����wf#ؾ	���?p`do�Ψ���Ӥ���֩GgWb��)ڱ�E�^;j�G-}<{�Q�(+��nSH�&@A�m3]lע�|�oe�o?�]8�_����a_J�oX��pngֵ�*�3](��3|N�|1jN�jh.D��OZ�8j^pA�5��*���X��J��;5�E�%s#���Cͻ��!('�O�Ʉ�G�V[֪�w�nBM�#Ry5S
B�BMh����<��ȋ�ϥ �����7����<{������˵��4���A�H�8��MXU���\��Ǎ'�O���Tq�َ��|�hGm�����b�T���9�8W�:����2�g�gM�Ӄe��;t�Bn�Y!���dٵ��
�r?�!:�'��ۀQ�I��v�\Hs�Q[ZsS�6���AW0$�r%�K��gSZ�N��5[����B!�����+ ��a9�o������._�F�3R%�K<{#C0�w�tޝ�9�Qd��+�����㖬^�'LЊ&8ap�@�}�!v��s��N7�	ПH����_q��7%�l뻉��P�%�t��N�o���&Ͷ��P�~��X$�#�����ŵ�O*Nf?�<���Z(d��`k����m�����pk����`��ǾV���`�2@��M��/{ApZ�'�_Юsp����?��%u7��=&9�>o�k��oL_�M9~$W�l��l��\�[��j�-^w2پL1�L���N_' W��p�����@9RlC���XASB}�qZQ��ћ}�:�Oߎ2+i�p��I�5�U~�M�]CC�'�t�U�^m*`�`yĥ�&��|�����%/y�H�͌�K�dѬ*�?�@ј�C���"'�t��=��o�(,u%5��NM�+����jelH]��3�nWM�?��}X����k�~:�:�;1���^؜��Y�W�4�z�����OMF�����Ǹ\6�0�oҦ_A�9�6�>�7O�zywWҊ]'�Cɔ%�2Aٖ�e�bZڗ6�������Z������Ҍ'h�oV~˖-|���O�$O�O�6�b����Yі*���x�Zr?�4kF#�C_�H͇���,9 �'9�p��B��v�c-b�����z,&��� ]F���k�$J2tp��{�9ԫ6�Q�k�Xx��	��&��(#�����0�{2��I���h���m޼zm8�2�yB4�R�^w��p1 2I.[��t���B;,	�%�V��נ8ݏfJS��sk�b�5�זL��N��N���<��5:�Q���#�o�*���O�������E�4��R6�b���� Ŋ��LF<3_�"�En�y��N.蒳j��D�B>aǭ��ѧc���r�l��&�&��Ϋ~�t�-�u�D~��-zx��d�֖��|��b�O�����H�=�7�JS]����m��.�?��{"+��骥A����Q~���AI��lrC���0�يi)�,98N�3V��wj'R�۳�Z�泖i��C5c.�0�Z�K��%�|<���&��vّ�/���,ݾ��Z�l �(]T�Q[+�|���#D<ig;�&[A���s�D��AKY-�Y;8�3j�~xT7Z���bw5(��LM����a�E܀�qBX�j`�Ie��s������G�V����QQbm���U�R�ûgZ�d8����?��Ϳ�	p0�[�s}\R@�#�d>�Ov���T3y�4�'wVj���-����:���[F1[$<uR�L-aꖩ= ��=6�v��&B�Eɗ�	�qs6�Z�}Wu���}��o4e��d��,uN��!�4���ԕ�O�
�}
5�{zة�?���p�2���''FE]��i4@邗3�.�ȥ5Ƨχ)n2Ϧv�n���M���kG�������_ ����92�|�i��J_�Y�I֍���i�&�i�#�ʟA.̲�[����٢��]	LL�º��9j�(��c�d�d66F�|])���2`�(f�/��@[($�M6�y%Dv���m���t����~yPIӕྫྷ��C'������92��up��ѭ����xc6UX(0���iiո�bU~#���*��lw�9 ���j~����ȧ��~M2��A.p$�+���-��6��x����J���Ga�Q,[���(��֏w	7�o7����ȗ�n�^*~�e�F�I�Y��N�~_M�*&�z�ӍZ~�x]O�|=��eEv��������G8�.�3����\��o2�u�gga����[��t�dxG�e2�xꍎV/��;	֌�5���J뼀f4�VX\��vh�f�|�]�s�m^��[��ݚ�$3
�ύ��G�2�ğw �6�
Y��#�w*I����=Bo(��x�4�#B-�RN��%Pr~�&pr�P_�'�hq�|[�f��z��~�r��lF�	j�Ҹζ]T�1'����b&����xO(��5<Lgn����d��)y��bi��<Bpc�p��#Ns���̣� �R�Pğ5)�-h3]�z_#������;ny-0"Q����>��+�p�1�B(�����!�����6�zfO��~��N�|.�Bܙ�'��f�V꒢^>�c@|�R8wĂ���(��h6O�������kRb�z�F|�M���/�0�T�i�F�����7�!>�g֊�������W&�4
 E��9�ϰ�AJ�_6R�es�ƭ��y�D�T�.�I@�u����Ԓ�Κ�EN�&��%�>��C�E��3VY�c3�;�U#��~Mg[n���&�����1MDm%�.0�*	�}�#^ɯ��=)�0Z�,�ٰ��$Xia�"q��=�y�.t3�6ӄ��qR ?h��hB��|�SN9���e�s���S�����9$7�@�%��#��w��#��f��V��}���6��ԘA�����H��D��H%}�߰���hzK̎8Ud�1p�����T!2�6?0?W�~F	�6�)	,uM�gI[`��p�s�
i@S�{�%cط���@�F�43�T��C�K$f/��~M'�C����5d�� 	!#YI$��!������58�9��f�'�=Y{m�)�ګ�ܴ��V�c�-���83e9l���ie$!��]�����V9�c�ڞ���FŕP�����(��A���;/�',���.���� v�RsH��xO�s��-�R�
��m��|�_��<����f�*Q��Zy�Gj~*��ev۱�M<cp*�N׌ $"?�wv�/#�
V�%2�o\K��Kd߿���0���P��d��|���	�W�Gs(��Kw��	�������"�1������X��4[���/�hN�U�8�]T	��{0��N�: _�쿆k�������#��&1��o�Ӧf��PՄǠ��"�'�Ou��_�LR�iL8�M�و�������Ꝙ]La�\�M���W�>c��zL��l?Rx.�)/`	��چ����U;�K�h�F�LI��r(=��)K��c�g^�S�c�{
w�o�I�	��V\�
�����Ѽb�w|0])�����c����&>�aY��s+��c�LO�g���T�?��ڦ�;����Ţ��^��֒�R�{�Ͽ��ʐ��(z/��W�����\A`�I�Y��.Ch�X\����>�c�x�8��KB�����A󘃷"�L����l�-�bD��RB����D�����c3B���%F�͌���PM2�ؠ6z��(���ZÑs�{
Tʼ#��|+Fhgg9�����}	��ƍgr�|N��(�̌Zz[��e}����P]�Ob����>�m&����׮�m���}xq�ˎ.�����h�<��wZ8Y$KT�׮����K�nf���m`��H��t}si4�cwʿaGigZc��$���}D�ޏ"��]�Y���+�W	>����N�����J�����r�N�j_ y�&8������MNv��i�R��1n�F90�W
�]D{�۱_S	8�_:\r|�E`h��My�7ᙳ�5qB}�u��yLꟼ�h13T�n��bug*����C2�̪E#�pG=�~�b�/t�}^�^�0��Y�y9Q��j���#8�ޣ����|n���I�s{j�l�h2{T1nT��)|�� HX���;�!�DS�������'e�n�"������Ѷ,��k��1��rL��I�����Me�f�MՍ[JJm#=�K�a]���8I\b�K��K��H�N���߬���I��*�~��%lٯ���,�V��h܊fF~4*�H��OV�[��Т\~�l�|�g�]K�2?���	6Z��fHoEh�~�}��Ltu��������k!�T��H=4��Sp�O�h��P�!"̿��Z�^߽6΍v����x���?�T�/�c^.��� *}���Q�(�в�D���o���w���E�����M�W"*ߧ&!���0� �w�ۏ�zs|<􉽎	�ͥ�&K�,i�:�J�؏�V��f���cH�l��2+L�d�x�*Z�53*���خ��&�53�_[��>��?����g��ľ@kԖ���@�E1��^��߳ <SR�}�PԦ�KR��\/5���y�.�o;�M�bZє�?�99�TF>��3�B�"R���I��=�F��S߳;�gO���`P���hc�:�q�ǭqmd��#���ߟ�gK�W�?LU'՘��#8�u���S�q^�t��m�@_u�������*>�����&�J}OˬRq&>Z�*?V�0�u��Tn&�:;<9�7|�#\���LO�8v%d���+�5�Ҧ�G�.&%߷q�J�e�,������rdlǓ�oEEZ���.�� �����[�o���U-��}eð�	�LK�Mz��z��wy���"���rq����*2����/��|����7i�F���O0QDѫ�r�N�'�YƷ�
�"��=��
ŀ�����O2��Nh�&W=!���E�O��<Tŏ�>3|�~�C���7M7��F�����ˈ�S׷?dN����J�~�����f�o:�X�U2�(,������z��^8���)��XH�K� R_��Bf�ܾg��f���r��E�����ᅉ6����ّ'ti�~��ŷ��<�k(U®��N��h�	��Jv���� �>Z�gN�l�X����#Q�:b���5{6E��k����	��b֥7O���Joh%dO*�LP�Q!���₆�ӆ	ۭ.���^}��Ɏ��҈<:X�0�bǺ�F��D�O��FLz0�����B��&�����
���f��͜we�c�����
���˂@�����ow̐hv�y�(�R�"�o}�A\H$ؾ������D��K$���Z���f��gi��*,N���u�Hb��������v��*+�_ZD�z��5�_0�_���م�����s�G~�H�I��/�N:�\�cvH�E���R𢡊��FN	������@8����K8ReCg��[��@�ΎK�.�9i��B_�i�s���`x��kڃ*���-s׭y�d�ϻ"�E|�*_�(��s��Nq:E��w+[�c�Ԇ�o�=�k�V�������9�\#46&�Ry�4,��_���	4T�=C��MC7'p��̨L9u1R�*�y� ��8_0��p������I�P:��Ie>�;���}+�k(I��q��q<�T$&!�?ގ۲+����V���͒�e�G�Py�!��y��s���7U���~���h��4<M\�Mޓn^H'���3?�����:�▯ �9��6!�'�[�YƊ˾x�	������}%.D�(��6�J�ѿ/Z��q�Sa�\n�L�6;Y�;�r���A��3#x��4���Ky܃\|,��6vY��Y�ٛc�b#l�Q���\A�2A�kiZ��r�n>ޏ��ENb>^I���S�����PN�-�!����O-��L�BUt��R_}�I���Xνm�N�����O?�]�{��̱�'���9���>�M�u�|�t~��q�m4���o��eO��@�L�o�UN���Q�����X�]^:@s�{���'n3�K���ᓁ��%����w�k��iv��d���>~=�s�˘h��k?�LkZ�S�n���YH���;��_��٤���`:����xL.��c���k8x�[zh2Ya�Y=aOpK��j3!���>>ő���n��I�#�G%_���x��r�#���r�4B$cc����F6�Z�~����?��i|��5�l#�Vk��Re���L��;�^��yeR	���}��s��w��d�/��r$�U�-��	~��yH�]�S��D�T�������Im\��!���I�ɮ����̣q��f� ��9����y#�������vξ?�יU���ٓn&?n�@/��[/U0&⏼�v�cE1n�G�Jas�t8)��c}/�EG�u^x9�p�&�&��Z��Ԑ��IT�^��|5Yh�0��?X�׭�x�h`��W�F�g-ﮬ0РX�s?��<8�^���t�T�f	|�͟s�F�t~�ee**�t�Z���� �C5F�`�q�qtM�L5��{��/���
L�s�`�="�(����	mm����������;ᏟK�7i��D�_ڻ+�<>�j��� yWOƍ<8�`b^}a�[�̞�qR|wO(i����n�jf[��_���w�HŃ�^���4�.8y7����hZ;���ʏ�0������)j[�>�6�v�f�/��6�V�^�c%%�`�ߺykI���AZK�:�ȎP��ȬY5�O_�i����g�R�ST$~��l��̰n�}Q���^�,���o{)7���pܺ)�a���T8��ex�t��'�+��� �o*�<�z�Q�c�ȯ7�'1W�1�	�R
�9a~�p{E�v����u��7�\���n�I�<�3P&6�O;:��5	2�G���Ҭ���fj���?�g��Y`PQNe��-~�d��0VӶ=�&�b<�`�"t�aY2'�4�;k.�}��i}1�5W���7+	�˖���Ǽe	�33͊(���tNϚ�:�]��G�s��V�9CdN�B���Tb]��799lv5����M��a��V�I.�IN�v�2��s�%1�0h�<���e%e��}�;B�_��d��S,Yk_H���lT�qw�\��-�����FoMՍ����
P�CI;I�r:O�Y:�a,�:C+���Ԧg��S��GNƙA�q�{�>.����P?Հ��� 5�LgO\�^Ҳ�zl,bc�b�x����V����7����vv���G�-v���I�)oᇊ��W��i_���9^͏Ok�r�[jz�n|V��ߒ����8a��tX�jV�¦X��kN/N�o'�^�V�:���t�㰚���A��FW�M.ew�c�۬��8r�ȌbJ*�ۡ F�x
�A�J���Ə���S�~JP�yS�L#�9����l�ԁ�2{빯ے��Չ��#�>A�/�uX����0,?���p%�E�^��hu����7�/BI���{�Q:��ms1��t&�3+7�l��G&""�&�'̏a���=�(e
O7�7�z8��x��m�ϢS�8�54~�5�[�g�t���G
&s2��ڡe��=���v��C)� ܘ���y�)F¸��4w
cm���d��>�������i�l{�M��j��|�!D�]P�=Z����_�Y�[������}��u�OL���v���އ6b��!r4�����ޕ:ϓ'*r��z������_ob��&yY"��,��p�6I�q��ސ��&ZZ���Rv���!�zj�?St��E�`[�qU60�� UH��ѸS�E��dR~�˵w�%C�v��҉���~u�D0��(�:�E��@� �۰��@��I�]�hA-�t����-�0��s�Ħr%s��_Bw��G�<��A���)� ���;$.Y���~x�|ɊQ�iՋf.h�g�f+V�F�vо�Y�#��{�&��r��k��OP�_^L���n�I��Ѹ�������Dmv/�[1�3���k4����&�
��v,j�巼Mf���9�us1O�ʆ"J��b�$�-�������f��V�5ݎE�h��nJQքĴM���z}��s1u�00޸	>��Z+�A*�	�5�a�t j7\���,�!� ����Y=����sJ �e���$�c���\�&�ꛐWk(Q?���}5�����f`����L�Y�M�E�Y��c~5�!�K�j�x�rH.�<���4�_Po3w����1�˾�_�������y�T��Î8~}:VL�Y3��[H����u�z,a��.�����".������(#�ڞ������o�j��:{�������d+�A�v����>Y	w�ʡ�9`Ǚ��L+�ĝ�p���*��Ô)[h����`,�5����3w+!&GR���dG�3���,��GX�DG��M��>����ۼ]������୼��}�R+m-�whDx+��k�+�	�H�a�+E�B�s��Ѱ$�wklE\�2��5A�/��su�G�f�)�q��� ׹k�e�+)*?��$�W7C>�-��ط/>��[^�1а���E)�E
f�}h,y
�~NXH\el4{����Z�J�&Z�2'��8Nqݯ�<la٬I��yNS�vY]�TY������D�����)y���H��^v/<��UN�`]��2\)B_M'#���  ��(�HA�mn�E3��2�ל�Ggc����&�t� }>��5�1�k�2j�v�I��mK�F;,�v�׬#Ams�S�f��)���oG�� �W^C[�@W���"rا��V~/���/��-�XJ�����w��]|=�V`0���9O#�
�y]�
.xv�{��7Z����%��SY�[w?×�9�	�~�y���y�P���끽 P5�G-tў��ǉ�����Xm��)\���L'���Ź�/v���-����(�𣓟��T
��H���A�R|>���^�R��U�(kl����t��Em���I�7��y\	���]�e��Bt6�̸�]��R�l��8I��MT���§��>�i+��#���c�8�g�j��O���ȅh���{ՒkH�>�׼�/�� �ل��6p���wyu6��:�LpCG
o}L�F7��N/��	��?x��}n�m���G�\�+�K2�u%R;73J.�a]d���vb�Ͱ��E)�/o�>S$�~
��h���Q�'Z�wNH�������
�g��6��4�y��<�i�jO.r���1Qu��>T�_��|�(�?�a�0�cF�¨S��΄�[�S��)��5� Dl��˿HP7�U�}���쉳��x8�>�3�:���Q�h�<�gK��t ���Yh�ő�eD��-�*��Wv�~����R#vB�];h/C�/��C"�{ΐ=>�����~&�e��&R��� �H�2Ц~�.F@���w�����)�Xo(�s?�b��)�5ߚ.�W�T��2,��2�_���#��5E���n�mre�y�2��c�.��$R=��+��ſ+G����d5�����M��ϥ���vhBn���~W���N�C�^�����QT�հp�?0�Q���&�i�t����{6�iajR���jA ���+1yE7%���ۊj��R���H�����ª>�:�.����E�sD'߳t�0���oZUn�����R
#���/��,�P���G�����J$BB��Ă�R��t|��܃�o��o�9qJ?��4�<8�+%�P'���-1~E��ѯ�#9��Dɻ�ԥf�]B�:�������`S9Xi��pE�o喻U�MVR��Q�� ?#-m M�%=i�t
Щ��bX>UNr։�����2H�G��w@X��|�$#{�ā`�X�*�]s��Ꜯ���c]������b��%�з�3���6�c�93�rY�3R�S����Ӏ)�Զ�����
^*y���-������$�D
E����;X|����k��޺�)�rw�
<<��t�ވl��}��F3�4�@}2#�5I����� H�q��pj���Ϟ ��zai/�!$TA������3Iz�	�.��f��ɖ9N��M��'dH���>�1Z��ֈG��+�>�[���N,,�E�m��ْ��Ri���|nv�MyT�'D�fn��+M�]S ]�s������z�怴f�G�J�p!��5ۼ&��gQa�H�s� ����@Y����GO������E�*.^mۼ^?8r������8�^�*��<���ߐ�
8��J�?�F*��JŞ���{�Ӄ�~ѐn����]�Q����ƻ�ϰsm��� �X�n.+;Q�DI|57f�j1z�v�֕�<�eD�(��$�;˪LM�u&�w+A�1n�IG��
%���ml��Q�H�����2��B�A5=hGq�
�s`QE[_�W� �+m�cy-�l��"Щ��N��Q������1y|��Z��L0�P{V�P���N��0�
g`p�У�\���Р�Ҋs�����䍡����J�s.���~�2xtwa��d�M�%L���wg�p�����Cu��G*_J�C�/�8BV�?��OĊd�4�9y[X�4����,�����B1_�:!;i�pB͓����B~��pY�Q%�;�dw���Z5ر��"��¿[5�E�P�YY�9W��R찂�T6Ŏ�'e�54l��<��Ŭ[�z�Z+H��:?���U���S"�ـ�HQe��p����j�G�M�ame��A�6�Ib�YH��H�V~�gH\�6}_�B�V��B+�m���.�	����xXn�H�����Pqh�"�47;?~��� ��y���ZH�׮��=;G1c��̀��Z����gh�����vrw�oY�8����&0H
{CuU�,��.}v�d;�$c��f�p�p��T��h��?���c�#'�/���	^��K�����(�o�Cs��W�*[���ȱ�tSbџ����fؓ��{Bgg��W�@�Yk��?��	�-�P�ߘK�KS�،�ڙ��$��84B�`���q>��\NҭX��eJ���V��;��^�그Օ�Ml9^��I��d,��2��\�Z%+�S�2S���K2�(S��������Y�v�|%L����1p�0`J����G��&���F�#X�L$/ـ$��0�5����\�ņ�B^m��zŅ>��3�����Z��J���K��}*�#Ťű�w-�[N�1Λ��.���r�Y�~R�2���bF�x2�=Xe��ScD;�o�B���؝no�"X9�Q@
=I��,�r�����?ϻۥ�_�������#�5��F��L��$H>��,j�Y���
���g��
��X��E�E�!XI�K��.��fA�޷�7.oz{��vY�A�D��( ��9�DM�Xڎ��k�tBJJ�P� O��b�tI�C���
�k}��u�؀v^~ϖ���I���x�u���{}�;C6���7���h"���űY՜�b��׬(���b,�.;W:E��g�H��>m�+`4fW5�ik��!V);�(�=�"����:bfo�,0҃ �D��Ix}�G4��}5�_�0��+e.��xxN;�d�?n��)���'��;��᝕�� �fs����5�� ����(`l
�����6lQ6;�����%����T��W��讲�ڧ�ЏZ���^C��Akѹ��P���۶|��jE����V���?�v#���Fb�� �]�>(���[ex�ķU�����T ,��`
�'+��4C�`�I�AS���x���q[h�(o�cŜ��W>��#l8��Wl��)8$�羀|�������,� �o���z�{ :��ҷ�Z�q�.F:*�<u��y�V�h�b��*춅S@��UE0x�	��C,���SYs�J�Si�����5�����u;��aFB(B���j�n%ROB����������O�VJ�?5D�$��p(�c)$Z�zU[���+��z�KJ��U7�ZDdN�*���`y��0ﳉ��w�(��Ӽ��e�AK��rq�.���
�}�'��5И�_����6�x�u�m��O(��.�.,�Y𵻆���������@��#�'��
����-#���`� �=�U-
6�F��	'h�^_t��sǬ��_3�� )cJpo��'.I����0'�T�T#���5�hmEir��AB��n���~2�eB�l=�C�|~���Yh(N.樍~�gꦕQb�ܗg�,leĤ�ß��ǐ˰����2"��y��5w*��T��	˵[�SR4p,m&��������s81��/t^*?���*T��H�z��m�Sh�gR-:qnpp4���so�d�T�����=�A]k4G\��\v!r����_�k[�RD(Ƣ\�E�o'��d"2���8�U��h��@d�[��0�œ66B5�B�0���ЏQp,ݪ�k��d.�_���wQ��(��{����kмAap*����e��a'J�e<���^�|"8xχ\}�0�VG;�l�0m@���KX~qm������63מ|.�d������O��#[�;���PD�8dc��,,I9�qް��t��7<��W.)>t�`��}|�Ps�9�[+�CE���rtR���6eQ�5	�L�O�f�&B�ɶ�_njá����֖u}�����fM�AL�ca�L�����٫Hጩ�˞��L�;V�\������<�ڝ$�Z��E������/�G	S���*�d8��%����� ��ȉ���\��Y5̯֚�[��~J6��L�\�D.��A�MC���6�hL@��<���1ڶ.O�t�W�N�I#�E9Fc�Rk���S����U��b =��C�U��u���(�	��}�ν���:Wo�p��y�7a~F� �P�:6��,���j~��j�b�� _/X?55L9��A#T���1(���EO"�_D���|�t��x�qŠtSܴb�C�&��v|�	s��j.L#,��-1X�JqR!���q���'F�'�}��8kjqơ�'�K5g�/�mӣ�34���uDy����{"K��Ç傐1�1�O�¿���3�a���XBzD�sW���U���q��yjg�T�I��Y�E���wWSn��j�G�kW��y",hb�r*��];.�h������f)����i��Ȉ���K�INwn��>n��3�bwb?<7���1c��|1n^k�a3��cWj�g7�֯�&x4W  �N�{��!h��s&�[+���?ULڻP�����缇���U'B^	���@�\��6����w��<A��9j�J.EE%���/����%c5j��;��R�75�E��0��s�sT�FFj�����WWu.'�&�S6$ �nQ^[^П����5E�����ds���䬢I3�Fq�B���xx�L�������Uf�^�j0���Bf���`��|c*���f^ܧ�9��ԢW�Y��G������q��Z�e9��;UKC��_�׮z� 0a�]U�����f��^5���m�q��a�D�D�S�w�2�E5�����d�U��b[���9�<����D�6N�x��5����W�6�[��N�HB|*�`t���ş$�
q���Ow��c�̂ȟ���s����ޔ�8>�%�������^���q��Kb�K��i�ao%���zw��P{����vgW�u���SL�/�~��=�:���)���M����~P���%�N���Q������ѩ��U���|ϧaA�k������S���^�ߕY5A���b>��/�Rc�"�<�;4e�������^���|� 9]�K�S�K�Ź�L�n�l+\��PZ$z �mS���t�
k��5���������J3;u�#~)��܅�<aS-:Ɇ?��_G;,jQq�#���\6z���#N�Z��Ӵ�9���#G-B!n+�gRC�)����C?*M� u���s\e|3�b?%�}��H���չ�u���̷�Ι��	��AD���&�x�)�Y�ve?le��������,[�Dx��A[�J`T��!{�g� >��\�(�t����1k�?�~�0��2?R��+�,���'*/��Y@@��Є��*���AK�[�/�'rN[,+�����c.���&��u�[��T�nV}�]�G�&Z��Hڏ��i�<�d9ͩMTLB�C�Xv��f3bP�4��ǈM��	����1�W���y��9�m�����7%���� ���Hv��7�ε#����|��_h*��OSю��ZJ���PRS>�]�u��pR��\;�gH񻙃��vh�D(d�}hOj�A�$�.�3���'V)��E�����FPZ���;�<*�ع�3�aj�`aCJ*���2КE�.@���GIK�	�`J��y&@b�"Z���8�6<����>1H�s�l�J#mj�g"�QE�j��>�Bh֝7t����Q ���wG�%���{p˳��i=Oʁ�J����7T�� 64���c|3�ɳMM@v�m�ɩx.\�99l�0:wjb���a�����O���cs]���i۩�!���NXw��5��0;ڈ����a�7j�iA��Rt�5��Yn��j��5��W�0cCꩦ�zy���[��0���+v��x6eў��+V$�y����/7�H_���gW�ma���	���5����w�3Xpw,�;A�������.���k=��>�?8��<��~o�]�	H}�
�ˏ��7$\m7�����4F$�1aj!��z,�b�����ے]���F�[x�X����W;Y'��%+�j����t�fû{(b(��� ?߅�������b�J��0�	S?i���Ų��_�&�zڡ��l|��	�ΣDA�SW/y;���O��گhnֲxO�6m��&��8��	�a��#����,�	����_/��6D�So���%= ��^ٮ�4^��hw�<���3�!���ܵ�|�����(@У�B�P�1�9�2�z&��clS$qR�p�&���@Q���XЅ	tv�A���w�S�>`���9�D3&#à�K$ģ�,���`�>����&��0V"1�K�l�&ԪH�e���\~c2����6U��_y+}�]+���A�pp��ZfTw�.��~u�u�(�ϙ�*Y��1�UO?l��ˍ�-�Z��\��'�����*p@~m��5}̽�g���JzA�X��d�W{���`�@!~ƅ�^%�p���x�o"H�M��ح�~��1�ߴovǓ�(B����8?�r�oQ_�Z��.��5�y��j���ǨI� R@�:� k>�7�ur3j�w��4{�j5�w3���@!�~���ǁ��N����.�!���9�펊m��F� �3H�@^M�1���"n�o%+�&��P�lmj3z��y��<.����Y�o�����X�m��-�e�n���_A{�z�*	Q�_�! r�=>��Ή>������Gq�c�_.�g?7W�e���,�&;��B�io��f���xwF]����e9X8N��du�p�.��!d�?3c6Y'��ꯥ[2��kz�O0pZO_�1�� 	fu�@I��(�Xs�o>�	(�X����Ν�Y�,�.�8�3!�+1m��׍�r�}�7��f�KjЯ%شG�v�	Q����P;^@ɨ����/2�&(8���E[ȑ�4x�.��O#۶Ip���Y%�z��&dE���`z��?f���E���9�<���P���dl�ḯ-۟�������$pZ����
���Ȝb1�����9�����9n2��nXM��֮���υ�r�!�v�R7�����f�����&+�gW�2��/p�߾��M�0C��G�R�H+9Ԅ�~�]RtAu�9�c]`�y�5�V6�ᡷ���#THz�I��(T�X5���D����|z��Q�v�]kW��D�maQo �~�J�f7�" 6^���Sʢ,�ǚ�{�~�<y.� �/ ����VZ�C!��3U���o9�`��k�-z��j��M���v_�G���q�'/ًe�ZL/0�3:���S�����t�ӬW�uE\T��W��R@�Zh/�{b��dY���e�ۚ�f��\n��[u�<�+����:kꨰ�:�G��N��FV��Ӓ6VX�5V{�
�x|�D_K ���� �_<�3�ͧV"]����w\SM��}H2Mq�b����̧u����Ӝ+�@~��LzYM� vj\U�y����[�:���3�����S�����`��:�A6�'�G�cuV�������1�������M��p��x���M��-��nխA7� ���L�H�vMw���N�jы�ɛ"V:�+��Ѻh�U�{s9����gI����2pD�c�2�ANLQa㞏���_�B�*������#	(�Ζ:e�[-�߮c���wv���8;xX��Y��=����{*���Յ9a-������C����ص�����z�378J�o˨��ۚ������o	�{���]~x�~�e�����D��9",s��3H7���e��y0/��*5g�|O�!tu�ȹ�j7������E=`U� Gq����.�G������t����g|j���͕EmwtL��Q��\�~�޺�n&Fi��Uux�'�5��,�Wq'���B��#�+pA�m��V��ͬ������SHA��V����8���P���!4������t2r��35�Db��g�9�zp>��,� �҉����{5�$�_H�qvo�~����Z"C���eL�xx�X6@,�{C�s`s����õ��iؓmf�A�y�*)�.0i�xoFW#X^��c��k!�������S>�e%��ĻF/�N����L�5��p�P���`��>[61(�����:P��c�� A�P8��9oE���A���n7em
Y�D&�/8�����.<�����!�deR6�����
���5��X�,C�!�P�]*�7�>)�|�ےa�M���բ!�o�[��y92C,M�&�ç\j�������i����>ΩK��������7.~�5��b�����a��<��o%j�K�}�1�D%�&���pt21ɹ@(B��:�"�Pm���
��uji�!��b�����ǘ��γ"�Dp�������S/�2��Ⱥ�W�GK�⹡N!��z[M�l��A�6X��?S/S� 6�9o��$-������>Wg�	�\P��b��Ano�>�,��p �$I?�?�[1y>��F�Q:�c5�����S�^��(xs��SPM��/�q1�sb���L�\�C l�@I�		��^��5�ɤ� C� ��?u)�nèS���3_2������ ��W�Nm���MЪ�`���\��d����]��Z>CE��`��ad��o
����&h4�Y���7
U��1?�̿+M�����U� @�3���?���'µ�:-�����n���%�X�mCf�0�k/�"�Y2�7_W�A앺��<��h��%�ǧ�[�vH4����-���%�������� ������Ĳ�zھ�g���M��&�����*yq�)�4 7�F������WO�Y��1	H�Nb�dǃ)?Cٽ)�R���B��O�u?r����`��䱛b���������6���vN��1G���P�?� LK�1
�	p/�AbX�,�Gǟ�l��9��<D=���ZJ*,���&��'���R,m2-kv�P�)H�xk z�-9���V�,]�6]��DM��F�}�Q�t��������!R�BF���'�,d�d��5s�����$͋~�r��Q��;�����	
|SF�w�����إ.{�+	����*v�	��F�ٝ���BPsCy���f!�wB{jw�Q���/���t�>��9	j �DY�AB=�I�_��q�Q5���h^�&g: Ew��Js�S���Ho���Ν����U'�f,Ԭ������:���)��7h`/:Q��e�����}��Ey�ғ���'��q��^�TP�Ly�������K�3YX��A���_�BW:�i�0�P���s�`u8����w޴��C>�����E�*�|�dr�WnejJOLi���t��zI&��*��o](N,<�a��2|X{"m�*k}82|;���@io�*�����~�/^G��}%\3�Z1?ܝC�!�d��J���8W-v@�����4Ph��xL�i:f�1XFZh����e�Ő�8rp�2������G�V��`!>Դ��E܋Ҵ��>���#�:��0LȔ@K�׈꽍U<>��I�p\��n� 'i��62f�A@��u�Y)'�9[9������i��V-ZK)������0�oD�`㭠�����ϳ憨L�d�K�-�|�@|�i�i͒*7��(;���fm�l��c�|�#<�B'�v�Q�R+��;[ו=��hĲ�)�ҎP1G��M�ݓ�����>G)�!�A�}I-C7��P�_�l�P!��1W�x�}fN+"{�j�Ҝ˺:ayW��|ś�i�Ɵ]��Iӂ]�lF�G��i�LZ��k��(ʐ5�p��a��Pz�&���b�������~�5M�h�}����X��	��B\o磫Rͧ|%n���I(;%��7���|���������~�w���R8McW����x7A�X�8[v�ynWJdǡ��<��F`p��R.Y]d��Xv�В߭GjA���~�&�ѡ�$�Ʋ!�_ɘ�c���P�	 ��RF�td@l��ʃ�K�,7�+���r�Js����W�0ID;;W]�'ymIR׍���G|A��I��[�ѵ�f#�JO�x��_ɷ�YŠ^cX�D�7c ����X�I[>Չ���	}�#��3xB�e�;r�Q�d�g(Xd��#�C��:V���3?�ThJ����R<el�?o��W����Z.� ?��I��mK�[<�г&{�?��sZ�{���e@0�p��`����㊜y慦^�d�Tn|�֘pCևG2F�I�ad��t[gf:2r�S����H�5�q?؄ư�r�K�A�'������wI����bQ>����U-�&M PY�@��cG���>�ǅ���r�#��DwHL�>qH��EJl�p�&Ȑ��lݚ��#��u�S����A��O^<��O���z�'�L��1e����j=ԚEu�� �����^�7虓{wV�:8�?f�uC"h��: �ۗ�M����C����7^ƕ$�Ņ���yJU�}?m_���Pk؇��vl�_�O��h�m�nI�u�?@��e�0_�Z��zf­�ܝ'���I�!��8\[z��ri�p�os �~ �5J5�dUУ�\��	4mj{�k޿.*�~�9�W[��C���.d��'�F��%�;­�?N�#&���������[�.��3��R��������\>����81Ǖ��.����ŲNg�Ǵ�RAB�7e 'C�A�F�4q���%ܹ���s36寨-!N
n��̥�SV^����_fg#�*��!�{Ͱ���O]�-rW:�8A�����-OIn�AI"��9�N�,A�<�+��{�k1h�,��!(�����Me�7�r8�Ĳ����ę�kgh�?���E͙hrv,e�5�nw �KbNB�A1=S���C䨝RR�$��xR�tzx��|�(1�i@���t���X�>�1���ϯ�Ԕ�����O\��v⟫�)�A9\��gF3�����9N�x���y���3j��~=�.j�&����d���ꚓ��[ַ}��o��I�)�1�x��D���0P<
/�9�u��c)����R�rZ��E��a�U������A�q.�"��*^��Ci¦L��Ǯ���0UՌ����t�?9ԥ�r)7�x��6��`����
��Ѵ�(��w	y��kQ&6��++3B���	��7��G�l�^�`���7�fz�C�ɎfJ�!x��c勻�Xr��u�������;�2޹e|���/�1�	����J��Q9��n�����(DN����VN�L>���T?��CrP�A��5���A��u#Ca7f�˶�,�a�8�Ռ�ABl�Bp�.�.��-*t��&N�N�$l:���!�c_����m�iy�W�A��ͣ4��#�G�ѷ]r��EҮ�,��:�;�����k��u>b^�DL�n�����{֩s�M*+q���{�my����xc.Id��f'��ؿ
Plc�}TD1z<��F�H�<6���/�<��uQYԤ0��4���"+�~�T�������\��!��N�Ҭs��<�#�w|�J�qc�����\r���D��w�Ш�wq�H��5����JŠ��G�d|s�B:���͈b.���E� j�k�8��S�N��q���oL�#�n\h���>?�Z̊ZpZ�a�VW�c�1	u�K��wp����2!�Rv,N�}="��;������n_���4���%���i�c�8�S9Y�²Ďa�)������A)�X6*��z��m�(C��OT�Iͥ��l��	Y���E�uik�����s�驪SKg&,`��,ʷwv�gvy�����;�C\?ȿzl�h�\���1��K�@/�`�����{}Si�����7��fԹ���G/�C�c|C�@���,eaD���/Ĺ�����ŗ�ӫ//���Z_��~!٩�<�C��j)�B�nF�Ix������b� WW9�y�7-E�P���2h^B ��'i�O�?bg�]�|^��1�=����*�濸�8w��9��r����|H�<�0���k�q�g�ot�uv�P)ɂ9��sIv����`K�N�F�ɤa�U��{�S~�5R��"&f����!��H�@ .څ_���R�:L��g�Tˡ��&�I|"�)� ��-3y gH�RЌ� ��U�����h��IN�?���ꡠ�-3:#��:gό L���>;�$ގl���c�3[#�@�l%Q�T�
AH!�-������W�U��BҌ	��D@`#������x0ٛb�_�G��Z�䝑mL�x����g�ǅ�	���7Zq�?�3L7���[��ӵ��-c���p1� ���)�dA)�Џ�Us�P�����D���^lM)�IO��\Ɠ�qt�\�m%G�6�����r�$]�L7��,ٞ5�����N�i���%,7�iMP�x�2��z^ �q����9d12�!����,�����i��/-f�v"x2=Y�Y{�����A��[�r5���,�ll�	?nA>cW������g����ۢ��;OP $d%�hw
8�sۢ_��<>�R	���G�з�wYle-��!6^�R�����=y���l��1^�F�	��y|��}D�*:|*?$�H<��)��#s;�|]-A|{+����4w�?�!݈v������Dt�zk�ǜ�M4��֒&GI� �fK�\�;��X#�*�gV;W����
� '8���Kk ��cd~ntV0�W�L$�܀%&XtԒ�n�����yX��c$<���ĿR4c��诀�z^
���y��Zk�ʣk*'�G5�f����E�
�ˋ`h'�T=q|��Bu�b����σk�C�F]���-!w�6Q��Dr��qW^'6��ѷ�<�D�67|"j���*aT��b\1b����s	�-�6��4�p���!�8��E�� u�ͮ������5�01��&�6w�l�1�x3�ď��D�2����S�{<
ٚ������םeذm�[����T�ͬs�����8�"�$rР��h\���4'�h���۞���y�N���x���	���|1Ϯ��0��E��9�n�(�[�Z��&bPW��i��D��'���o��}�Sf�EF�8I84b�)~&�P�r�Mnq���My>z�M�{þ��TX+�@B��]�Щ���E�K���p��z^!L3���5��Ôz_�`�Kmk��;QfUe3�����+����E��VK���qyi��=����-4�0��s��|yz����n���ߟ�r(.%*��y>���G����3�ebR0�R����=�'��5"�z��<]����X�p&��s�C���I�Ca�?TH\g�o�Q��\���S�<5��9�U�8<�Z�|�A���
�D��@���4̌.�c� ݀1G-#Vi6o��b=慖�?x�t��a��~�:Pa�|�W#�>#���v.��/<����I�����ȡ]䊝��r74gT|t�?��i�4m�(2T)���k����D���a�/D�ê���z�}<�������G��W�R+5���).$�!��K��	UL>ʶ�x���$�8"F�_�kH�9m!!��O��_F�8U!�^̷�(/�),��=c��v��7l��ǜn���fh*�ĝ�8f�F��M��,�	He�r���Urk����K�piQk���fu����K��C�����_�O �Kw�䍱��e�枩ob�B��B�U���H�h��{��dHVI��8��d��U
�wi�e�^���||�t�6e��4��D t۫`����E�	0���n�g���ˏ>��=�<��6��(��P��P����|��&�gFa�=3�z�/�ټ�S�^А��׷�uO���}�g~3�q_�!��t�{Q��f��.O�2��}�^��X3؇W��gVl��#)�k��r]m��r�d�C�C��0��j��6�g�
����KB��_��x�W�_y�_��Q�)yy���&�7|����$o�t�̞$�ǊT��>����(���y�Y^k�������ѽ� m(<��"G���g2hV�gG+�� ۰Ԯ��M��rк��Cu�m�4�B�Y5$����ݒp�����E��OS�v*�-�с�8�pv�z9�!���dkzx�c�W�o�m3ldL�����ۄ�؆�`��坆�ds�I��y�~⾲�J�5-�TS_���-����^�肋�=�Y��GJ��=rq�߶��P��M�E�j�1�7�k��]�þ<�E������1.�@ ����K�(�$<�#�ǘI�Tol��d]#xvҜ�1E���qᠢrR�z{�(AN��E���
���>�.8��$���N��V��O�b��l�~H�c�o�4p~UBj���Ĭ�0�5��u݌�VBtsԬ(j�'VM��x�����ʻћ��4����	Ԏ6ks?%�X�Gd$�.gh�f�-����M���i���N!&v���m�ԲS/�|1[�7����g����@}	2�C��V�3�]ۉ��0}M��t�
JT�A;YA>�엸�H�5��w��)� �Hf��/�182��nh��'N�^_�l�J�ԴUx���e�ʘ������޼�;�~?���D%�B�i��"}�U�����%N*�^Za�A�"�g�}�;T�&��Q4��i�E��kq 4�p�>��?�NN��K��ch/	�����v���IT �v6D=aU�s��8=Q�g8��p�c>5o�r��z�|S!a�����!�� VyLjq���b�m_���.��!�@ѽ�"-SJ��� 4P1�._��_�Ճ��̂�Y�^>�0������d�m���o��M��XDΙ����s)�(3U���lG����#�Rᶎs ��!6c n�T�>���+�>�Un�����g u>}��'2���*��f N��Jym[I�j]������q�5ާ��*@ T��yks�s�;o��\��� �6�4�E��SV�R
}L[��c�^&d���]co���.В��$�������j�Wh_�K�s�br!
N�#��e��Qw��7Q˸Q�^[6�;�p�������xR�E��`Ƃ���մ)*>�q㗕0H�9��vv�L�'tfŘ��t�0.� ~����($�?���,�NRx���X�#�([�u,o������%�f��2���=��y��	��"$�w��5�!�
�냢F왉LfqU�ɢ�� �F��']jV�OS7����m���X���9_�^�v��֦L��(,�@s�N���8�+�i�9�C��&�}Qt3=\����s��Z�JT|X���j9�[[%/]��:������x�6sd��[�,��0��YR1z��n�!��m;��	X��͟[b�,�鵝&~�	�{�|�M�������}p
Y����x�bՊ7sD�<���KR/��uE�Z���ԳE�T�0e��",�Yv�Z\�` ���:�1�����ɀ�|�38jL��G�S���y�}�+9��h�0�,�l�1Z���k�5N��(�b�֌��/�l�	�K��0��krf���Ѩ�˅k��7Z:z'���F��%X,� xpe~���j�B`Yv�_��^���^�j����J��5K�qt@��.�0_��C�����z���iz�����ؘ'�>�$1J	!���wXa��J�Rn�0CO�,��2��buE���Dz_ɱpd��>e����G?�7�U�	c�8y�m�u����:��f�8s���n#
���ɚ �A��N��PE���z�~>�tٞ�'�4.�1=�Ko���f�KjX�@N���㯎x4��sI���ڋ���ZHH�U`�����7ǵ�aS���Ӄ.���ߠn� ��`-���vv�a��&� ��:A	�L�z2����;�ť����^�����;�!��!�`A������;D!^ۓ�P؃3�#��.�x���Pz�xu���lp��L�rڷ�
�q?iEK�;��/W��A`�APPZ����Hl@�ZH�"Sߞ�1�sɄhNr��c�F՗���r������@GPEK�m7^(����ݾЋxCXsy���P�ʐ~~Kd�%C��?AT8ޡ�z�7��v��!ɖ��|)�%�Bx���Yp��	hi�6��6^!�����I�f�{ސP�FKk|�/z�P٩�26%��f���|���;ĸ�.�*��j�c�� �U@{+��h�t1Q.*zF�ᾗ$����R�$��j���B=� 0�쇦���p;5*��6�߹r� ן`��]�ML"a5���aDٖQ�L�e�'�����H�������=y��e|̕��~f���~�ˇ�W<s1�2HN�!K�7�.at�Āy<��˔�oq�� 3[��<5��?�R�ؽz�7^���H�����:{�SsF;��&e�X�h�h������f �l�j��Z�������QR�H��Zu�YM��D�Q�׫��@�>��
�"��m��O���,��|M?s>�"qK��� rG&�˾_��$�zʅ��XW��#��ՄgK��_������{�n�J�L~�f-G1�9|�Pk8q=��{om�9�D�Q����DT`�v}	q�����KZ_#�4��!�O�0-�~�in��<a
<v��"�o�%�_���O¾E"��%�z�vz���s����ޒr]j�b�3k�z2";{ ��e�q\Ty�(�5Nj^�a|�P�ݨ_��f�u��ǃ�9V����]�g0��"s�]�N����*�vLX>H��(o�`����w�0��Z��uf��HVіx�?�Lܕ��=kl���F�j�?�B�,ae��7ǖM������C���vꀘ{<	���QKc'g���8ejO4� 	a^��"��	�`f�螉#�HXq��Kh��KkC{V,� -x'_�;����>~�f�Ý�=�$v��j���ty��c`ʀ���DeQo�T����"��O5����.��a�o-//����7�\�}"9Ӈ��S=��ER�(<'��䷲{`�ҏ���r�����~� 8^��op�מ�Mequ���s�β��������"�-��$̈r�ԅ���t�8� "��$�<
��Wb�T+�Q�b�1`]�᳠�2y����h�u� ����ys��	[�2̚~o��s��˿�W����M��3,SSaDq�zkj^e���V�K˕�E�f�(�1Q} H"��!� [߉j�d3�<Գ�W+T�Ɠ+[Z_n*��	�8�]��ӥv�<O��N�aiO`g76ysţS�?C񎴖��9kK��a�����s��1	��O��&
	��Q��D~�VH֌�'���+�yR�@\����4��8X�3O���N������l9׿H�s��Y��Ā��֒�j>L�Sg��h��<r��d?���Cz.~z����=� zDl<�ϗY����wߎ�poo�@��n\IE��X��w%�|J夵����{s}<�iHg���TT��� �l����\�e坪��{�W-���K�/��N2������qDXtʯ55FAHO�h�:<��x�K�����Wl�p%���O ��M�����p^�����y��|�a�^&� ."�ÿ�����=B{EU"k�iqPϢ�g��d�5�^��<R}����}`�v�ک����$�q� c�M�E�鰎�q{��z}"Fb�m�W��\َP��MQ�~�^s{����?���R��$|s���)a�b�p���K}�gi]���1r�x�ʟ�L���}?�;;�p��B�[��H��&�c1��2w�:��/�?��7%����hp�O�.^|��h��NU
��u�G�3�U�m}�e	QVa
Iܦ!R0�Zi����D��@f{jШB�#�#�++)߾
=ǐ9�-�\CE��s�L��܏�@���𓉺�0d�Ri��/^��~�R$��q�QŒx��hK(^V�vK��`ysPI�%�L�0��Y#$1��b��=�
26QÄq}	T͓u���.��t��e�555�^Ӏ!P�+:����M���TO��0ތQ]+9�!��:n����	��1~
��8��б�n3������5;^�4�6�0|,�^��´䱚�)D��+�Rcy8�1�X�$��Q4`X�Z	:M��a�"r���e$fG�Du��Yx�T,"e��!7�a@��.�4E�8����/�&|��,�P?\���g�k/S��͙$x�b�n�V���4���'/��8�~���@ `�������|ng���s�����m�ʲ�J�}���D�c��"��G����
���Z��|f�L���R}%�}L��N��t-I��k��c�ǆ 9�S�����@ˡ�sK;)eg��(3�X��)I�*�r9̓)���[�]l���fѦϛH���h>}����ʔ�(���Ⱦ�]K�(���D�!�E\:s^��?o�n�9q�y�3�+w���l-�v��,n�E~��s�v���۟ٸ�.�i�I�8rӉ�f����������=8���l��Dx�px��u�\{����P��j���c��MA���^����0z��FLpA�ay\_ U�����e�?��Y���v�W���{��[6�_R�5����Ha�8���(�h��5�I����k��t���t��>����B}�v-9I��٬���Ӵ�[0�܌�"��J,�7�Vośc����~����Ā�R}��u���ፃ��Y��@/����A�������B�Ṣ�Z2) '�<s���y��JE\`�'S�J�3��4c�hnd��d���t�X�����$�����u��v0Nd��wW�1Z�vvq� ��ש>X�μ��h;9�ю-\�u�92�+��Ե!�@r� ]�ߢ#��bZ��&�������/�*IF��;��2���=g8tmll~S|Z2�}�F.j⬈�ɚ$f{*f�tN�J>��M|���J�:\���������k��WA�V�\�s����K��㜹P��i������Ij�-7�K؎��r�Ak������w�$�mP�y�ܐ�n�Ŵ������?�����Z�2���������-*��Ȇ��Z��J�Gg�e 7�[�t\����~�?W��A[#�/��^���=�x�1Yeg��xk����2f����x�V�\�81�X�}ܓɴ,�qL?vM_�z��ifl�tu���b�a�l��	גj�|����
\ ��.��m�J
��ԟ�3�e7E��N���r����q8������~����[*�RL�D��FH�	Y����˜(����@��F�B���N�ʵ�`U��.�'VB��6Ω�����]`�P^�����+m̔�Q�'n���u�S�Sm�=Tkjj:1x0`��+��u'�V�젫rƫ��N4��\؂,��|t�I�E�U�y�FO0�#�3�c�-%�Ԃ�߮Ka�!'=['�C7VCsf"��9�h���(^%��_�����HL����Q�-UF؄N����L�ܻ:���.�c���x-�<�81t�.��j��n���g�eb�0q,T�7п|q�h��l.�t���d$�}�G�~u�c��@��>��|2B�7��Չ*-}���ݔ�o ���,���]ڄ�"�X�Q�$�`y���Õy����:@z5�eCݕj#B���a�����z�T>-ɖ¶l�n�0ҙND�����Tr/�M���4~4Y�M�m8Q,,�1��"��m#�]����,��l)�.1���G�}�v��;+��?M����LO�u}+s�Y�!H_���f��Z�U�xD�:�3o��������vpe��`�/���w���&	�2!i{eFKY��
�\$p�/�Z�%�ϿB�'�"�_��V=2-�L�XL+�޼_;y>*����jrq��H2J>��M=E�MD-��-
 ��=y������e�?�w�K�����{��䯴!ӭA��J���@e���(Pmʌk�b!�i�EZ?�n1�+i�[;��>��O=VX�4����	��E?~�9�9'��\Y��,khgR���5�AW�=�1Բ�N�aC����*_�e�[%�:c���������K5[V��<v\a<���i�����,����j����+�/Z��T�5��p�Ϗ�)K2�cL?͑�C72��B�frvs�/�]���� ���SV���;�������f�,��	E���y��E(ϒ���m�uO��-���K��ȒnV	��7�9�ҳ�6��	k���(ޖ�J�mH�
���J��Ϭ/��'��?k�,ꑜ�`����Xv��ij܄Uv��AJ��bHҡ�86MD�"u[dΌ���D��E�j���aT�>rI�jK���)�NՕ;l�b�V�#�$�Ώ;L1�F{�R�&?���6��J�S)x�z�MӤ��+�F4�9��n&J�-��]���ƛ���AC����]���Y=#��P�	�4���.D�_�)P���kX�6 F��v� U�6�cv��_B��ޟC�"���(�T�,Y�k_��\<x��������;��\h�h��PGg��G��-���l)��ܟۘ��j!>���z8i\�/��Mb>
>�)���Igk��;^'�8P���^�|�:�Ȃ��~05��V���8�i6����<@(y��b�"o�#M�ٙ�X�fT�5Q��*���J������ٺ��3�֝��"�z�<n�ƈhi-z'��- ��7]q���>�X��U��ə�mi�cS���Q�V���g�d*Kpo����m���i���
�ι��[��mc��y���.V"%ۻ3~�D�߶/�_���"�=O��fT��=�+k�íZ����#sH����^p�^Q�p��b.��!��H �j�a_�̐�!�籿�t1ҡ~<;h8�Җ����^kmDʊ�,N�#��=��8e� 'tI�=�FH�ᤞ֊��A��=a���aB�����0���8e�u��I5�,5���s{4���k����;O�3��x��
����|��H���c��-��(����G����C��p�Ը�	���|x`�V{N,lm5}_��|r�	\tX�PS5�̴I�^��\��vz*�qõ��'ƅ�6~�5xwO��a�a<&���ʀ����L��$���M*��>e��G�'h"���I9Io��f{�\|V��iE�в�{���̴0LTN�������ye��;��u�:]۽�'ǋ�8�o(y�
��fJ�FḡMk��
%U�`I�����U��c�	C�OfE�s�"���ȔrM��=4��g�H����\'N��)a?��g-�8G��$���2��PޅBJ��yI�6S\I0��D�;��jIi�:��g�7��=e��-,C��q�+�9���F?�� P��^�@��H��TdI�+�
'{����{�VB��AK䅒��cLI�K��*���yd�,4u��U		}�J(�4�i��rR�G(iI��!O붞"�#+ߪ�m:�ƭ������<�2I?���.��)|ў��D8���P��?k���"�iL�Mņ� 2�\\郘���Ƶ%�1�k�M�bKE�)�|Q��2.n1�aw9��l{NO׻ۍ�W��м"y�,0����Fw� r�|��[�!O7�u��՜�(?�cV#�b\|9�[vg3�;�λ�J�Z��Z�)��Rt�l�cUT웮ˏo���RlYֆ�yo�jS"��}[97�fA��@�(#Z������Χi�:��� �z�K�h��פ�:.�8�rs��X�s!^7ѳ^�4P����@W?�G�i3�l��D�)��~�����[0/�,8���fiR���D����\���C�ɓ�]RQ��"�@`U(�P����)I>�5y�G�_����H����Zၢ8�>
���
I�u���
+���Q�,j�*�N�An��/K��n#��Q����	'�Xۘ�A�@�c2��  �͋w�H��+���g�+�H�^T�H޵��#V.�w���6�[b�9�%�̤4�ޚ����Ä%>PH�Kir��bZ�ZG���*����IeO��a\�I�4��ݦ.	.�#�ո�hp�"r�zr�Hlӑ��b����SѨ5K���?����x[e�f��$�M퉾 [.��OWEse��"w���c3��N��	I�q��h��1}���V�ǙP�����v���F�gw���"�g�,�5��_�X�q���.�?���8�+�zϋ�dy\�c�w��+��]��.X���$�AKv�e&��rT�l[�sp���ֽ��3jp�>��7�*�T������\r�v6{��S��8���h�������vseվ��*��k9ySт�S�j)q���⫂���q-n(���Bq��%h�"ťP\���b�w����}�=g�\䂋0�}�Y��w�Y���)(m����1bjA���5��II%�Eld�J)z@����̰�����W#�R-��Z�PW�y(<=k]�S�0>��|a�Y8��Ϧ�ty���vl>V��c���4��]�nN�N�9�Μ�{���P��f���iv�1�� /�&<zPI�N����Ra�q}M��2����l��6�\uXܯ�7�F� 
6�!ڭ��
��#>{�bp�7�|���I��Ub�ě&�_e�v��|;)����򃐲�=���eq��u�nċR�z���w|_Ŕ�(��@�.�?������o(��`���z�8��z{cF�϶?�)�Z3�8xJߧ���w{n)�����vcŏgo2���5������1�� ���́}�e]3���}����V�>b�ٓR���� a�����-�l��<��'��`Ď�ƻOuZn��Q:K��C�=gE� ck+�7)t��ZIK�\�y�gO����{i����8�	G�ߢab����w�I�����fH�:�b����41�"�
���_�w�4�'Q�~�L�������{�?�lN�G�UK��wCU���b�A��/#��X�x����y�A�`���tۤh�LᏥ�[c�
w_LX�}�lUK��̊V��)����$�G�%I�7�G==���|�`q���[f@��=pE<�.�M��z�@EL?�����yŏ�d_�s���`��x��f�����J�8!nG��{���,m���?�h�����"l����)��Jkߙk�@��ښ`j$�����Q*�7�#~*��(���	9��_G��j��O�Ve��0��"�(�`�5|�3*4J����I�J���c��^���U��}x����B_u:�2~��-K~���o���1���;�l�>��r�$B�9�H����|��A4��l4�@7�����x*/p���)��'��9,��m!���q��������QK���V�kJ���EL��7������0�������X4_��|������&����!G�K%��t��7���ɶ� B��p������/#A"L���e�+�ッl*��P���jOD�\�o$��P��c��0c(z�-�S�����mT(�KZAzi��}���<�Q�[D�o�"�aL.sA�4���'���Q�bP ��;���-�))y�u���4��?ԇK�Hj�7�t$�N]����'�K1rb�QbU=Yx>�]H.�&/(�	[;f(�l�Mya!!�Y������xV�X'/��1�H�J8�����wA���e*���Q��f�b�?�9,}�w�|/�2��N#��q�ǃ��D�^*e]I��- -sHr��N�0����g���p#���n�p5O*����}��[t��8<��1j=���<�:��τ\��V�毝�E�� ����1�(㳜��^����v�T���I>�a�eآ���⯢�%�.x��{w��+�J������/��k_���6��D$jX�-��H�����4)kڂ)�zzzn0$��+���t�:�yg�\+={N`�#� P�r��Z�(����̼_�q��ֵ���bn�§{$�d1��~�kN.?*e�5���M���>M+������'v�� ��i䓙O������l{�?vt�ñz8)0��{�����l�|�H��S����Ü
 b��6J���E%��6�����	�|���M0y�xTe�=j�h�'։f�B,���ϐ�wu���)<�j��Uö��:=�ϣQ�oz##��cB9�m��ׁ� ��������z�(�v�Y��~9j[�92�xZkU�[e����L;	l|�o�YdXsעSH$��&}V�^T�}@1-��Fah-��k<��?
��V����L�X���ޕ�{*Uґ��NH� ow�0�t�y�H���p�_}G�r,DI.B�d1t�2{���=��$\�j��%^��uϰ#!B)2��AޖG �\����KŹ�����Qs��y���a�%��H�k����Nx(G��6Ï�C���4���'��%�������s�-ܧ5vZ��*��(>�����Ȉэ$�d���93aL�E����"0�!د�����K����$\1�G��ύ,�����^#�� ,S1,K��	����z��B(D��)�*�T�"����6 ��3^5�T?h9R˭��H�r_o��r�R �:���Q(m�V!�;BjU,�@td�:ak�]-����O#z��������.<[�S�����^QKY�x�$�Qc���]�^�^���P��ˆ��c!���ޞ�	�#��-��K��	t�F�5rV�i,L�ʋ��N�^$@�����6�r���$����ɭ0�"�~���� ��H����BB�D�R��b�A��o���v��R~�sk�|2�.Z�Y 6�G�p\*��k���'�@��oCc��I�7C8."��BG5gp����>������&,���J�I->#���S�K��O~�J/Ye�5���_��������H�{�-�!���;�9}QV�X�͖�fՠp���~�u�)ѹkS#nd��S?�ƛ��y�y�| P��� �����lN�6v]�K�#������o�!��呕�A�.vR ]�LA4 ��"G���J#�ߏ��p>��7��>>��XI���YH���f��tx�z�V�im���������L���y���y���Z{;AO���Jk�U��
`�h#a���'�E�r ^s	����w��Ǘ?����aƋ��ql�[�(���Y��)�T��;���ڥ�༑�E����e���M9{��%�bz����������1Z�i|Z�쪌����s�������t\�*S���ذ�$���T��Xjh'���7�Rܕ��-���Z)� X�4��%�������B�Ӑ��/�g��(��NRL�@q���B�Z.�%�K�tl�S�Ҿ�h�D�}���$/-rt��A^�f:Ñ�=��n=����Z��b��%�+�~gݲ�#��W�s�C�<t�#�1��P�\�� ����J�M�K� 6,!p�#j=w{�����ڲg�сO�f?��%Eo�C�~Zr��ח`�T�t!��<i�����T)^�5;�c�U�mbo�]��c,ŵ���"/���/������|?v����*�C7a�3�q�pk�n>R�>G��"e;z�{��Grataɬ��6R�<��A��1Ŀ��0t	�I��Fd��(�DƱ��g�Z��K�c",zB�o�I��aY�1�X�t�J��+n�"����	=�55��%��}j����L'�EzH�'�o�P�J��<�	�G�V�i��>s(�U~�h�j!I-���B�f�7,���Sܹa|��c���XD��1-��Y��>��h�|?ů�!�H
	Z�%ܮ3~���QK���n���q�b���XT�����m�&��Db@��_@L�\U��:�f$�{A��9NlMb�P��_Ɠ�>�\�|�	��U9ԔX_[��$z�c
0~��k�H�������'�\��^X�2?��h�����tW�Q�����y���N?zB�S�tF�0E���¨?��Aʹ:�w�c*/��>�gz�:aࢹ��J���&$	����u�I01�w,�!�~
�
Q��X}�U��ƚ��b�=0|P�+�I��{`h����}u�?���I�����h΋#��B�
ٿ��q`1S�r���5gi�f\ng=��O,�4�&*�DbGg@)1�mO,��}�`i;Cp�����o��	\j_ a��P����1����oဠȻ��Y������\���-�m8kXR	Бk��!�X�L���?d�`���ԯݦ~���h�E=oAw������-s��Z���,�f��?/���>��٭����	F�Q*Ø;K%ײL�����y�kC��@=�_YC�pb����(��{b8@MwCa0�����u��#�W�S�b6��|��E���}�w͔��b5*���R��^��M�"��` #�2���,b�����=�~���ؔra�\�m[� ,
�6'�IO����*�����(�:�A�=�M0]�&��-����c	 '׾dz4�dx��	b(�-�̠Fs����O�x ��TE�/5�SL��>:�X?a7��{�}�� ���2�X��ck�ޜ��P�b�* �cA�Ń~޷H%��ͨY X3g����"��8(�Xq[�����`�\��m�4�i��BG�N鄤��A��:w����k?���|�,V��#�l�2�&��K@F22	u�Z_M�4 �x��!��}�(�'���ڪ]m�6s�e����K�.��?F���&|ZAy�:�S�0��X���=%y N�"�f���R2C���W���o@:~գ���a�����Km�\JO��TG�ֳ��Z�)pޕ��]Ra�̇Bu�w:������b��A���_)�~Ќ���l��Io���Sh���{����n) �x������{�X3*�O�(�J���`b�d:D ��E�l
}��d��qzw�1������e��R�ͮA�Ǝ��o�n�#�-}s� =J��ŉ�G�¤�_��F���DU����j�#�΅@��'��+}�<a2��֚���s��!���9B*���V��v���zV�D�S��v��qJVSP�c逵�@3�y'�ɼU�:��œ�2]'�#>��|��uQ��y�����b9�+ڿ��JYm闏R�M�, �理:
�n�i�
b��q-M�j�#U��￵h�aХ��[��=[���f�@�(1y��x��B2n�U�deC�cl�o7�Z�"�&�L��, �;�~��O�Ƶ;�I`�=}^'O�q��O/�J8x���������B)�60e�0��#��8�C�g��7���8�H5�l��i��$�[ ��^��'�Ն_u`�2c��
!ϴ��@Xl���`��D� 	ռ�̢eF�OCr� �|���o�'eJF���8�>oP���K}�[�Lm�����/���o0�'�Y ]0q���v�|�<�;��z��ׁN)s���F*���J�d\�����$d�+g���?7����ѹh��Zno������C|�� �y��l��v�VⳎC�.W+N�s5�Aj�v'.=�6;��.�樍�%�m�`豶�vd�>Ix��1��}��l$�r�?�~�:N?1�o�q4O=9'm�pjy̰y��
��=9Nv�e��@&�K��ߘ��	"���@���	��g� � V;�ü�F}�cԂ�^A(�.��'��.��	I1�#A0 ����}�e%�D��]�h�H�`M��������+-��2������-�\ˠ֎vw�pi�����$�i	 C����'$����R䵋yBv$ .!o	�yd���Ѹ�v�t��.*Z��o.������bG?�cE����x[-��V��g�		Ǜ�ͯL��5������)�
�!�.�
��ǎ�_*���4� iz2��į�ˬ�_#D��=Wshu�1�NG��J��!���e]��y����:G���7�/Zb=8����ͨ=A�	ͦφKĮ�{L��-��&���].G$�����m�g`J�B`��-����Do�� ��r^�7$8��J�`#Be=ќȕ��q�����Q���Q���C�ۘ�����5��raZ���(� �Вٓ�}_�S��u�t-��߿�c��V��恭w�C�H�!Rd��~�Y���#�]�޻Ź1O��X��>�C�7��/[)\����k��||��j7��V�uњ��o��bT�yM�l����XY��k�+\�l�o"d��a&�A.�LE�.��lg��"|�H�D��N�5��d	z�r~8�UL$�,;6at.j�J&���I��R�̍|��FV�]��A->�;��J�����+&}Gظ*� ��n�����3/���|��2m2��)��ƙg5
���7|k�B�Mb�?�':fr{�u+���μeR��փf�6J��߸�? �X�a�n��bZ*º�}����!�mc�:���f^-�=9R��aIO	*Ð���噅�7]2��� ��ͧ�O&_�6�Ѻ��`VQצ����4����.�2�?F'. x��F��ޏ|Bfbը��b���X�S��_Z+�B��U/[*��g���E�aI0���~`;	���y������Ri�/�e�#),Y:NX���k�3Ÿm���&^"���1�۾��ȏ�~ aD�i���(Z~��O���`W�Zvv�Mlh���ܪ�!#P�֘p����R���=�w�4X�����9�ƕ?�Okb��F��Y F�ϗH�;��@]�D1�~/�0�x=^��yMYv�1�81���܄�|s@�l&�\$29
89h�E��n{4[��#�0�s?� �4���}��NO,�\�wBU����b�!&/��d�0��ڈ�B�� .�5��|����m���-m'�#P�o�tj��;0+�^ �-Q|�׆�b��hd~��6v�/��%����j�����A���+��O�0�?��-�!GO\�4�C�����D~�J�e"~�aoO���E�����&MH6�n��jez�[�ߎ�f9���P����룅�.UUc).�2��m��c=4�M~nK�s����i��=�$�|)�c�k�~����ڹ��	Y�M% ��|�䚹N1JfH;��X	�ޏ^4]͓R?�z�l0� �t2𦶓�:�,v�m< �ji�2�XbH�p.mi6��N@�h���Cm_��F@{����	2��X8x�zÉ�h���sl{O���d^����-l�Y��0���:�v���b�ڮ�:�UBu�!���X2��o�4"�_P(~3ӹ+���a @���`-`#���9Q��X{���q]@C��j���������|l@�h���_{N�کB����B�c{\���J��v�=�}D��o,S������_�P�/�aՆ��J�v���YL�}Y��Dօ4�D	�<��B�yM����)��d0q��\���;�Q#@(.C�}��߱5!tst��!p�S�΁m��ý
ϴI�[Ë���^�q��BB������t�]/?�޺��yM]m�on=�H0S�|�O�����f�Ci耄�@��R"����G؄������e��D��HY۱Y�:�)MWbC�i�94�K�`�fZ�&��5?~l��䈸2_K	i�y̙�ނ+����f�N��2���N)��������V��|Q�-A�>�?��np�����s�Pw�,GүS����#�*{��,Oa}��8�D'�3mN�-c�H����|1�ߧ��$R�t�D�I�7���o��I>۝h�mAs�'����!�:��a$8�>��4��R4��B�� ��y�4�<֧�M"X�
�qJ�MÈ��LD2@fH\Y�b���꭭��ޓ[�혎պ3f0�j��Up��Q/4���7�U�Л�d�ߌ�Y}�.�Ka���9Ef?���-���ގ�&�I��K:�4_��p��
���ceCoR�����Y��h��� p
������������Ș 1��?��`*�X��n��B��d���;��!w��6�˿(�-�ҙm�V�@~t����ѴW�ᇏ�Y8p�b��Q@����n�M���\9��.���TI�k"�W�� ����5�iV��hQن%����A�T������[�Y��ڛ�}�D��dG��\�65#dg)Ɩ�#(�u��Ey�2�^9yyҘ��-d����'��Ε��0e�ףY�ga䳟�޹��l�C�io,C���t 0V����,�`�u�<����HUNl�����k�iK�KnJn���r���ͯ�G�ب?
��#cT������s�pռM6���i�,Y����ӗ�WV@�-[N��Ge*AI�-��K\��T�F�mS�N�N)�{$�?���Ey�j�!"MZ���`hϮz2��u�ԓ�D��"Uzw��u��_8������;R�s��Pi���Y]�*E6~��:F�aC;��Ycw�y��OO�$v�y43b���m��	���"�rX��"�7FB@+]�R�b~w;W'�Pɿ�����-���Z�\�t�l�hJ����閆���|v_S����������ch*��>?�h���s/+�]����h�&����EB]�JQ�ơ��H8��؅d�p�`F�sޒ���Gy������a$��-$V�3��<~��3E%� 	��0�iU�S�&�`��*и�� �@v=�K��Te��(λNP1����3z���_�?>A��] 'C�%��ѡ>��Jk�8]�TcNçH2%��Ha�T]<L��D8��^��G`ᥐO�U���ӎ�U<"�����	
e7|W@�w�j����<��F�S�o�Ҩ��Ԛϣ����:�5ԀY�??9�O~�zw9<]d2y_��y;A��5A�U��w���Cb:��kY�N�=c���5W����Y*id��v�s��)��X(��iF���w�]hi�90��vI��ͳ�(�VLQM�.o�.g@;Bn���. �9�N�3�Y|?���Ii[S�_4�KORDDd�7����$''��[���"ɨk����R�L_�:�p5�
�i�=�����L��b#�
�y�%�]�_! ���tݔm����jc�Oˋ�OQ�V���>�ASJ����/�����|��=�O��׭�k,`��T�L]@�d�m�C��^AX���JK_3��@Y�<[�&7�� �+4+���
�����W�s��N_�Ĕ�)ǭ�w�JߠC��Kp�L��C�������{F1-��6p3��݁~�Χ���
��jU8WCW�����i�7��34�Ӥ��`�-X4��Sv=)�FfX��Ϩ���9J��wܳ؀��C	~k���wq[�/=Dys�l�>�8qN&(���)QxW g�j��*0&�s���*'��y�ig>LXe��(?�ap���L��ݕz����Ht�'e�I�-������L���yE��M0g��4���u������r�Ǹ�W��rgԯ^Eq�\���z����Q;k��H�L��.��������(����l����$Ї.+g(�h;�EP}UE�+���vzj	�ޏ??Mm������Y�-�;�қ�vP��ء��@ǿP�Ho�{�j�������LA����I�����Vȣ�: ��x�f�8k��,�т����FʅY1�5��D�ƪ!�k7��u[mꋺEC�L�U1�|j�ױmYX^�:6�����TBmw����N���\�gB#��2thQ��S��*��Țɉ�O�՟��IYu���׾0E[�!���J@"c� �!7��W��AE���2:��p����	?ǝ6,�7O#\��d�Y�"�េx�b��	�ᄲ�TUǈ���@Q���6)�����#�����J�)�����2���xT;uB�A�詇����>0�$���f8��-P�=uvd�ƍ<��J��{@yR6$����h�8��\��{�s��4c�[��;<�{8�&�jA@�2<��zZt�F���zk�G`���-���?����J�-���N	�����&����q�(t�^@�g�$�B�wcW/0���{|޻�ַ~�]�!���i�=Q�"���cf���e�ü
���}�D���.m����ثֽk���9ɞ��40�Ž��@'�Rʓ� ���,O�^}������Q>H��M䯕����k�H�kn��zp�5�~'*�[{Urǝ���c$��q��N����ܝ�������}-}*n����'7���o���}O�i��v��}��2�Qr;{���i��"�}��>�;��}��e�7X���W�D��˟���Xk��w~��6���B�!ȸ^$o�`3iN��M)N�y��ӗU'l���.��C�#�
!@�P��'�xmD�`���:q.���Zn_�FGȺ���|����7 m��ɝ��A ���J2�8��忲���gN_�aѴx�z}��!��N�L�1�[�~磱��-��}X��=���s��)\��G�U�C��e����@0�Ϳ���;3ǘ#��J�g7(`��)��>�S)y��.!�&�/��	���6u��K4t������x�3o�C5��{y��"��)�0 ��x�.�GbK]F`����6~��'���5Q�g[r��rG����Iq$�w&HB̉9��7��3eM��((�ۧ�y���������t?:��I �a`s���{�8x��8܁�-8��K4-V����`���f#��?�J���[.Ɍ�,�Hb��6r�6�4��$k����&_�Fτ�K�	����{�N爢�����>���3����Q5��8l�x��X���7td&ze��AX,��C�E�X}-c�*:��ز|����zwmѹY�}[z�٩��7T�&�zD�{S��p%4����v���~���J������VDN��;0�r#TC枮���ȅ����/OD=�J�0�eJ�V,���x�u.��Y&�����ϱ%���u:v�)Khi��k�T�r�0K���!t0�����f=C��c��_�D۰%hP&�RsrM_	���t���y>b_r	��v=�l/��Y5V��,�]����[�0�O.�v-�*m��sZ�2�7�Da�a�n����D���l9䚪OE����U�� �$'�@��|�k�C��#�W����"
%=�eg�L��|!�+E��ͯ=���x[��z�;v�z0V�B�s�� ����L:��]RG��L -��ٖzL�� �z
�i����M	"`��nk���%���b�4*�f���	�h�sϟ���,AE�E9��-���Wn���۰Їf#SW����k|v�7�=F��;h�4��č�|l�k����3¼�ҭm�����c���&T��r=�f/Y"�,-,	ɉ��<��(�7����NH-0��-�v�nM�-�
��0�S�Z��4LȖ��괐�Q�Qv&(��b����w`y�UBV75C��܃됒��qwז�+bS�S��$���Q�5��ȩ��N�UY����������z08a�;a�t��w�F�$B�K�|����Ʈ�J��8hȢ��5��S��)�(<>�����_�G��*�����>�tGғ[��m�0J�hm����E��?,v� 3��O2Dgwk= ��J9Γ�%�h��d
��T��y�X�SOʈ�5�A�e�ϕL��|i�RT~����<N��ȷ��ea~\M��~���^����}T'\��6v�!	����@vx%~YG�<�p�՗=�=��돭������eN�Q�W����1{��|XO�(�K�&�΅9<��U��4s��t:�{�@}ԉށ� �GXM��^�~S�.��0X�<��n���z���$:$3޿�ӓ�4"EFoM����!�9๷'~[t?�v����p��k��sr�����z�y����������#����\j��))4򼅣�].~���u�´��r�%(�����N�r��T;���,�`f�JV�6��ˀE?v�	߈����A��q�ҍf�vr��{+&Z��ƅ��+\�u�6���b��8/�m����i��������EM��	@����S�����bЛ-�J��7�^����RH�H�Y�&���^�)O�N�9�W��W��LuYV�0��ƴv:xg�k�Y�ז�N��J95Tw6��72�M�]����N0w|����S�����i';�Ŷ�;P~4^"^EN���=�E\��t	���>���!��wB���*y��%�1���{��;��1-E��F�� �����#j���Eҥ}0�gUqQ�X��Y3�?�׹�?�&M����D�<ߺ�h�����À�>T�-Z��%�}���*X�nP�����ۘ�O����4:M��D��X{$'l����@�mY�Lu�I�����B!֕�&�䇎^ eB�^�X��vR�_�}/�Qj�;R�����>�!s?7���6#��̡IZ����2����t�ypA��K�ڵ�����
�&$R��V	l�;MsjP�����/���*�:���9_�`�E���Kg������&���7�y��r$�{-�N�4����a�m��3�Ґ�>ǈ�fD�s}|o�ɛ��{�%����fhH�xH��{��Q�ǿ���z͉��8��������ss�n��}�#3N���y5fZ��,�兰'/s�5�!Ik]�H�'����qiEt���?����yא�L��8�[��:��_
ڂ�����K��F|B���Ð��׵��׫ѥ�#�)/~- b�?����e�֪^~c&��O�U;��'�7n���Ae�ւĞF��0u�k��6ݺ�;lJd�� h"aJ��m�����}�]����
x��~����w���FTXK獛'��3���a|a�(�� ��J�V)�W�i�T�z�j���e$熲7�8��۵yS�JZ�zdU$&q�g�&�̈�j�؛�Ly>��~� �Qg��\�=�́��L��:nͼU����m/�e6�1�F��K%�fY2��Y<)��Ff���Q`Y���&"�<��UU t��;�T�S�%�C�e��9�_7`$��X��ށ��Ž��TLx��	)s��^�߿�y�B������g�e{��u齲�Dih�����+�x��21	�k�]�O�2��u�����7>��\A�Z!e��{yJG�5��%-Z��6�r�o����Jb�����4��,���SVZ$��6�I�Q�p*5آ��oL��+�nc�k�<��_ފ.��t��S�M�$�������,E������es�S� �e?ɋ�Mp����3*sYމ�º$�C���I|�S���/��$����[I �r���C�_;�BΦP}cv�<|dO9h��,>�X)�� ���vP�ؤ#����ĸ�c�'���K@����o�A#��q�T��K���yxy����%��,�����+I�bo�<|��hPU{���6Q��0M
x�߬�L���bԮ)nL��*u��Ǉ�Q�Y����o��8���v�;�a�L� ha��C�|�8����h��ɵ�<.�d,OͫA˱�<͎�T�N�KUx���ӄI���'?�K1Ok��u�����#x���L��^��oܙ�V��[.��|������bLi�.|�n�g��i���W��e��!���Z����p~&������������_�`g����X&`���k�g�
��C������tF\�Q���u�p~G�+��W6�Mo{�q�������+�O�1&�7����).Q>
;	_#�2v�L�H�\c�4�{h�_ڂ���ݺ���9���0�j`GyY��ֹ��
)Z)F|Sp���U�ȔP���/��9{ݩ�6^y��[~�j(*����L��P��T�MJ�5���[;�@�G,�%�ΡK`�)'�A%���6��lL<�����B�*��h�:�/1��\�u�;��8ǗŦ��$!�ɷ�ͻq��Wܼ�5o�߭R�H�Ă��W ����HX�e��Ug&Yw[����9)p�/�]z��LJֱ7co����S��9��5��{;.����H�<`鹩a5��v4w�yDn�I���t���1��0�B��(�V��O�;�F�]��r�r�>�z�z��}~������M�ωcي��lD�@�}�� J�*��;l��e����Wx2N�4��[/O�s]B����˽������!����
5܅�~�5FRyh���q�s�/��-,����	dy�J���ߴ:`N��P=kX����:���c3�*AԆ�� �eDy���Ӑ׍�e� @�V*��f�@�W��7	_i"��v�?hΒc��R�b�V��D���F�i�n��_�c�x����>���SNB}�_{/i�p[��f~�S%��7�ɲIbٺ����օU����v��Q�-��3!�/�#}�e>�R�,�TG�����tW�ֽ
Q���Q$ ��#�`!�F�(�I67[�YL�W��Xy�8?�>�+�+u�����t�#���4#v�?�� ���եLs�V�6� I���E��,O2�&_�#CI����n U���e����-�(�_� ��w��7�Ч�Xt�up�n����e���dKvߓ[���u���(��uW5�
M�����Y6�s���nS�w�|���W�}'�1ƨB[��8��)	�]���T,;yI�,jAu-�m
�+3��Na4{�]��\�ke\	⸟]
��ͫ�_�\�a��l��W�S��v��a'�V���� t>�d��^�.��3WO�W�o��hG�Q�5���+��u�[�U�
G����c������~�,0I�b�ϲ�#��w�8�v�S@3�U~������O?ݒ����i1��T����B����1hm��oK=�x��z���|"4��x�I�SC3���#��Ês1��OhT�{����}OwN���&ע���ƋAW+�5�ynx؆�f��<(��_��I�Ǉ��v7D�6�|.#��9'm�N��kF�y�α���/�}�)�[K�d��u�؝=:��Ж��[�ZU������R�Vh�xR�튵�Y����=euTW��ab�,%�T4����5װ���#�~����"�7�;�����_^�ja�ɯ8�:���H����7N�n���R�g=<����1 @m�M��R�B�#�9�a>��ǩ�Y�G>��>1tnc��-l�{t�p���|�Q�&z�N�dҀ��e+d���#�z'\BL��h�tE����95JJ��]V����q��o���'���gO����L(�[?����:_+��3	��/?v�	�1m�g*�<]�O,�X_�;�BŘw�L�W_��2�j�hW�����	.�����e�j�ݰ%�a�Q�̑f��S5����b ���َ�.�1=wz6���Ա�|\;��j�#W̌�K}�#��̵���vM�7�;*��P�a>���40���E�G��	�Gnѡ-#��Sz4�iq��ϹkQ�P2�k3ߺ`�D8F�6q�&�����&�����X����x]�ۄ��U��ZZ��?ʻ�r��umcD ��\�@6wO���$M���bb�8(�/g�&�꼆�@����F�؍��ՠ1�]�U]���d�a];x��3K����i��p�;�.f��q[�����oB�b��$$��kaG�`����v�O~���T�#�9�
�ӊnS�0s7��ơ"���'C�p4q�{�S�m���f��>�.�h�.T�d��;�v���������C��a�@�Z@��tؒs�X�A3}��R��/bS���ô���*O��?�w�J��]�Go<���6�����J��ogRI�;N�l��6�F1���x�@��c�Uו�XC#D1�x�M?W���V�edmT�U7&�����{=ўB!9�%�C�~���)�=�ȡk�1>z�n$�p�`��g]�MG��lc9��EF�*�������-*�&��; p@KEtO$R��3��^)}�q?�@���@���3~�[ȟ��ŧ�X^b1DҸ��r�U��-Oߎ���g�l� ��Z�������~��3>Z>A/��?��*�f�s�D�X�9�.��2^�:uc3�������T]>69��WDGE������3�u<����#��W���G��7��}P��R��I�P���S�#C+���������#�j0�ۀ��[���o��c�'x�8��#�Q���v�ۆhI1$1'��8�K��}����~vA�����W�"J6��_�Q�n�q��HJ#���n$��:��^����CIv�&�m�2XRNh��J'AZz���8�U<eILTx�}_�ː�ѡ�c��AQ..ZY�7��r��uccp�˗���Uy��@$�o�0 �[?h����LO4��v7z���p����N�D�Q���GD���W�qb���C��9�ex�-'�k+�q������d�ul�*��Uڴ�O�IW��5�{(���3�|�{�]�D�4'~8�,�ǒr�	�ݣJ����fNC[[	֟�����yɢ0�d�uShzn�WD�f����wl���[	*g�?�81N��b��&"���`�t0����>2���tc�l�5T-�6�/<R��X��_�㡵(���j3ު6_��ũ	��?V�	����-3½'p�y�������>�~�g'�����Xg��\�� ���;��dl��~�P��0e��ub;�L/;���oj+����n�"�|��U(��хqǖ�z!�
�;tQɷA�}ɛ��mj�$�� !p��U��п��ȧ��+}�ܱ��*��)˫)vK��MgG�tm�-���%xpܒ@pw�6Xp4�{p�n���A�������A��t�]�jݵ��6	\��(��]zz>�	�d��l]�1M2[ۓ�!���4����'�H(z�jÓOmֆZZk�,%���ZS�[r���z�
�X
�v�{/_�~
wo �3�CL%1��p0����c�}{$��j��$�^��W�Y�����p`��!�n��)VQ�z�6p�i�4�x��WA����	�b�5yn�F����SrĹu]`q��Er��Fo�#L��^󎙑\mt��o�T��[��_��,'�KTp�آ�9�p��?��D^��l	d8,�����O5�I�<��M����qr�e�����]!��;���F�lӊy��L�>��s��lfL䣧��oV��@s�s�P��9�׉r�L3�q�~��ǔ�\�L��s[����µ��y���f_�j
&�v��uö������n��fM�xn,�2(��NyIz���?�ЁK�)��Gr�QLVе�1ӢXt��Ɖ�[�~ѣ�2�!5}K�L'W�!%��)C~���wA�C�� �Q��X���-����}��y����:;űcI�Jc
�=`�ލj]v�o?p���F�5�Z�I&�F��]"���Z�F?������a�P��
x�-�����w��v�|��Lk��ɘ��V��2AmV�Ө<{�x,Z��S�C]l�?zq)�M���=�a�2���03-�΃~����X������J�lՔy��2����X0X���d[1�����&UV
��dK	��8�O������n}U���Cgotj��zjDx�S���Y[��w�{<"����mkOp�p��}7[�(0�Ͽae��
��Ӹ@M-��[R����%���}�#[M#i�jc"=?�F��XVĺ8J���L.+qy�"1��y������ʉ�?���"(  �ܯ�F�{*%-Oإ���+�𚘐����<Z���^N��{��.�a����w��nĨ�O7n����������b��]+�<�^�t�76kHK�d�3�+�V|}Gy ��V���"t�o���=������,C�w#��ݻEL,卵\��d��lQ��&?	�kK�K\�eR���:4��݈z�W�����{0��g��;} f֬K�;j�A�����n y�d��������x�d�,M,q��86�0E�T��,0%-EE�>��$���E��;�a���ΕN2��xFo�7��H���&���,WK��ws_��X�׃��Ձf6��^.0�4�r���d��*��:X���3��.7���dF����ޮ����\�3���e������^=XH��h6�X�~tJ�x������ƎL�0T����?��e�Y�*h�vS�����5##��p@^�E_��3Ғ��W�T�������h�r���mx�H|0v�L9�
����wQ�_`�����I��#�$��۵�# �j�8:�x�Q�����]����G�9Ud&5%)RZ�ϴuML,+�GC
V��"�I��Ş�������]������y��xΈ�/�.pY�M0�m��^
�߭"E�m��x��NTDH_=ת�R\B���h@N�w�;v�=^�m3<j�(�v8�����Z#i%gDl�F���\ �$ro�8u��Z��0F��J�'���<YtqJp(@<#���.5+L}f�BiL�sr�Q����wS.�ң�S�DG�`(&�[�*��d1 ��y-t�DN���N�_��{>������z,r����^�FzNG+�O;���4��=�{ЦȌR�XW�E/�����~u����9����3�EN-Jy�s���fW^A-ܩEt�L�9�mL{y������j����\��-Q�����M^��.v'�g��̸VNC�X������	��L�>�z�\\vh���I�b�6�f��h���SP<�����E�����^�����j�p)���9c���:���.>����k\����}����\O�L��1�)�ɯ��0�e@Υ�$ݗ>���J��ȸ�=�����ꛑ�0�F�w��:a�lC��z��+�s���؊22Ǘ��ꂞ����ө�`6�wˏ�3�}�p�=M�{/�ɉ��e'd��Uvdh䪕�饏�y�E���V�
l��a.�J��ì{^��C�ơ�;fIƊK��� �٥�&���@�����t��P�S��b����(ٍ=��	�^5�-5�|8�5Ė���g(ף�hem�с\�-��z/�j��R��^������}���-��G����<��~'��Q	)C��q�������3⍄
A�j%��
��m"�еO�k'c�-��P4�7�ȵ-�⾜=Me#~yьK�]�ywt�{{��5�����A,����p����,�mh;B�Oe:UNv��HK�6=��f��z�^�`F����㯴�I�-59���k[+����UL���0η�!��(?�`�z�L��	T�Y�rQ#����W���������j$Rpbu��(' *Y�-	/�B�]0���*���e���]���FF�/��h]t�����Ql}	BqDpLR�Ľ7y�A��5�_rs�F� �ϝ	⻃\�C�A�׍p;��⋐�/_���#0�t�`�3�j����ԉ~�%O��Ww��~�8L���V3�W��>j�įϿ���BԶ��[-	�ם��@� ��6�n��#��]�߹Q�[M^�'ْ%}a���
z��s�a4��G6�A&�� ��-�J,��[�����8�{)�$h�W=�3����z�G�����%�=r��nk��T�ߦ��! {߫^S��ȉ%m��u��_�����n�qVRum��c�~�Z�R
5�(�]��`��y=�����c�m�m���t<�JkAo�]����PH��^�����w��kz�$k���PP�b=�/ظ�C�H 	^Od���;�-o3�y%Ye�Ebv���DW������(a&Z�T������� ��pv��+����aa�A�.����"]K���D}^!V�h����^C�4�M�2���4�=��t��a�&��x��K��/x���&d��w�k�=f��Y8/�BV��>��e�Ã�jؤ._�_^�����让���!�R�zЭƬ
�^�����r9�KLIL���Q�~VmJ �\�����mq��)�"����u�e�W�w
�z"R0? �F������Fʤ%�b������#<f��V�Q`�esBZ^N�k?x٤������y3I�l?��ɉ�p��/˕����=
�Kʤʫ4v�0s���M�t{څ��������//ZB3=�Π��#E9��R���!��͜uq���*Ic�`�G6�b����y�k���d��@[��<�~B�� ��&�楝ؐ3�D}v/���S����ZX���������sO���"�h�mC�$�h$6�0���S���ͬ��������pԵ��,���`�:���ꀱ��kx��5�P�x;AQ��,�#��e�7�y>%J���1��g����ZZ$���[���9��޿Tvy����'~�5����jH5	L�G��*a���+J�:�Xs�f��zzlm��]W����(ǎN��~�����TW�ID �x�HU�{Zt�fªgo�����.�]��4���;ĸ��������6�� ˙�Ҋ��t	4��������M�ɶ��\.{��J�j׼ې������&�;�*���"`IHr�EF�=㸉�O�m�����<]|]jO޿�D�rf������'��.h	d_u���7޿Ai����0�O!�@����0aƝ[��WZ�=s�G����nm��*	1�|�1��6P�aŚS���k�D�/��|���/���2�j�7w�,r��e�i�*��d1<\>m>�.,cӆｎD36���O�w��m�p�BM������Ԛ�@��'O����6@������'�G1#�q_�����;jƏ�P�A�roڔ���$��>�`綱+Y�����4r�|>x�f�<J��c�
:�5�|m�~�X 
�^�Ng��q6δ�Hעh׃$h'	��,i��*v�0��o%��P���JM�E�Fsƥ��bX��3f��#(0�;�N{?9�����"8�A��lǀ`
���#\����`S���4g"���U~��'��w'��q�͍�Wol���p�H�eY����m��+�^'V�n�F=��ž1t���l���3���9��k��bR����[���z{	3D��aWF�rE@�B�'��H�P6E]	���R�䍳fC�fX��E�E�V"x&ۃ����tV=��%1�Vcc��r.�3t��g{�����Ř�p̣�ɇy��eg�m�e)�,��a�6��b7�
��ݰ�qN�]"9ý�p��
�ta�%�?�A�&��
jy���'v�{s���I�t�&�����o��~I�}.�}��)�JK��J�X[Bm}
[!�(�V��E�:��F�>�SOj�;�n��-��sP\*�N�"\����Sd�%�ۗo~2
v=��N�2��Z����O���U�}�m�f,�aK�r��k��9��n�:�§��ws.!�ZrP�#�3�%%H�]�[:-zm:��䈽|u�����f��?@�N�\�k:�In�����Bt٥#?b�=W��~�2Rb>;$�4��䂹�L_Դw��N'�|y���0殧vi|�aKA���`�ܔZ"����~�Z�e�0ۮ���÷E-g/����R�Z� ="�Y>��,�\�Сx��� � YY]:7=F����@��,��o@��'���=����`�+&���1����&���܌]Ǌ�N'\�-����6�.�IO`��O�{|j��,�\w�+4��n�{�T��Vn����
�KgL�r+�'Y���A���r�@l5r��Wy�[����,ǒ���I�������=~�i���Q��P�q_�	�[�)R�#A\y�j������ߢ`�Ӱ<-�op7��?�+�h��	��m?�I"��H���wz���Z�qʊ����0���cG����#}ʂn��G.[�ɧ���5�ӹU�z�}���M^a�a
l\��r<����EM��;�iNH����7O�}U��ˋ�
e�IxV��-b���4LL���q��n�./{V�@��6��E��sĵM�P2��~ ��0�I4���G`S�k}�{#��_�q�]���@����E�Xbɼ�"���/��M����-���~�����|Δ�P�������
5P^)B;_��~�:A��G������"NsAG)�����k��'1
�X�p-h�v�1������!+�H�C�Kn�j��v6/�h����TH�ʯ��9��D�{��EuL�z�����o����J|�"����c�So���~�է��zV�#��f��d^�M�jE����겈�hUj�:2_�g�u�[L������F�ؓ*�-.��\J|��4?�u��S��tA�2y���F��@�e�i��o��Z����nM���sN��AA6��d]k���G�HxA�I4�{���NBFu�q����'}|p������]"&�>Հ�'�2����M���VhQݹfʧ(���%_��Z���١l}3�	d�I�9��w�C6���(!^��I��c�Qb0�MT\����9]�No�N-��ZQ�������+��Fhk��\*!B�Ue���!'��
Kd���gQ����&'ins��������$������o��Y_��rP�?��`S�I��ej���;��j��7	�&���	�\�� iΏ�´�d�U�A �S].aW��0^���w?� �<�ݵ�������II��e!9M����i��Ȧx�Sr��љ �����1:�B���{̢���~<l��	��~�>c�Ӎ)�;��O��(<*t�!h��v�x�'+�n�d_,����j���CB��t���"Z����T0�c� B��؜R�{?�A�L|���ƒ6����]׵�[jrn�2l�y�B=e��mH��U�S��T�N� ��N_�������c��{�@ t!�`t���P�����!�q��ԯ�ʲ>9��,{ŧJ٧F��.u��[�׾�g�P|��`y��G��=.?t�ӁSqr���S��
�<m�=�y�M �h��ߣ�Wwx,@��7>.�C�k�^�!j�)G�s-c��]��z8S���nр{��=/�܃�]t�����U%�;�m�8���zӔ�#�R�����M �\�v�zU�.�ٜd��rW���M�y2�|s��^�|��k�BLp1��?��^��o�(\���1Aj$�����1���A�$|�v�!V�h^��O�j��yL�}<6��|&�8��|�[�Ҧ�ۡ+3���s@ֽ5Z�򖭠/����*3�l������`d�In���&2	vj9�_�z �;�e���������q@F��np�A�`�L��:F���p,���53��68����/E��`�����A��M-�8V6�5~� ��2Ҷ��7l�ib�	ç�<�OΈ0oI��ӝ7��cnhn�#CsoQ���>�7��r�n�8�䳉��6-���F$I��n�bE{5�;���{�ETՑxr��_Eܘp�Td����Ś��z����j� 2��pG�C��[}m���:���?)��'��J2��fc����Og�@�v�|�׆ǳ�}��*�-ۜ�~���v��FjV�~�dI��<�ט�1���� ESG'�{G_���+>���6)��O�(�#������5�qt׫�jm������%��������h���|��������7���_v�Qp0IW4Qb�5�QQx:<{u�(���fS�'O� �
)��HEM ��\�_�I�P�A}+��I�(տ$��To[>0�Y�T7�np*��䚞e�/�%��>crol����A��4��A�#5�3}���Y*��`Z�D|�%��(22�_�ӽLVD��)�\3?����GʑZȅ:Xt$3�zTl57���gv���;��Y��QP`w�i��������]��:����T"uT��*z�J70|��`9��ϩM��k��ɷ�:��߷��(�˥��3�t*e�]	�l�فd��)!�q�a���&�d��~Z���}7�H�(�m��I�z\�3���t*q4��p�����=j����䂡ʦX'M��6��R�#����� �������r029�ښʞ�p���Z��@#������W��oS�\!=�[���B�Gw&0������˞E��:�y� J�m֒v_>>.�ܲ�սz�.��ok�fY�s��S��/��z�;��J�צ?9L�67:���df�p!�=����R���gˌ�c�=���s�GZN��B&�����k�P9@���go,���?(���RP���6�l��<ps�_�������tԑJ�u��eX�̮�����|�w�-_�?)|\0u�a��b�3��ȢN���P�]�k��O=�?k0;N���4����	ADa0��ր��Q�m�t�2�?$����M��,Ʃ�N��*x�g3�8V9�'<ԕ?�(0a�:QE;d�6�g���5{{�C��`�ל�a}Rb��_I�e�qʚ�m�߭	�Gt��#���u���}�1l2�����\/GM�������-�K� �iX��]s���؁��b���tȿ4��m��o����zR�[g�G��[�\��q�-Bq֏��(~X&
��$E��c�k��y��W�2K~j�3 T�Z§3u�Ҡ�J��Ɠ��v��gr�#I�"��ki��~:	 <)����T����n�/ܠkl�� \���Ap�ݣ+!?�2�,c��u������	��dtD�ϮT��&&�8�%�"��^�
�!|�m6��*��3��+��r&S9���w���H���'Mv�&+�L�� �����.���G_i;�`}�M�(A�@&�F�h��C����x}|o�w�4����r��5l�+��B��7��\���(�����_~L�`Gݺ�#�"���V���9��3=���waKa�F8�k�����>K`��$��r7�L�iON~�e�8��`�Oi:kF�F�d�Vǆ����"��h��l�H�|+�zK�ß�#�i��ɜ�{��<a۪�>e�m��w����UC�O<q�I>*�A�&��������µ���q�k@~K�����]�r��*��풊���-?���r:��� �n(+�97�g+�e����5)�c�aR�Eׂ�]<I5�.��e��Jv������Ot�P'�Y�-	.`���3�^����53��Ě&h�V��,V��Ӽ��]��9m�m��<���8k�>���������i*#����"��+�zC��K.X��>�Y��9��������6��h]R�W�(��y��涒�膧��ZF�f���]�o�k�gB(�_�ab�����m`џiM�*Z�e�2�³��jbTk�a'7�������q�8ۆǑ�
ޘ.��Nz�J�۲��y��z�i����^=+��T�6�։<���*R�v�0��c���zN��'S#ӂ�$5�7�c-u�n8n-M0J��UV�z�r���y�*��.�ݲ
��qQ�ԣ����sT���>Z
��؉6��۽ĝ?�+�Ы����z-���6n<��u����d�qY���s4W>�5�	�S�,��'6��u0�6K<b��M8�UT`Ai���ډV�G�N��w1��i:�[
ʷ��e����'�y����E�shp�A�������V��M��W:<�$�zA���Kی]m؀g"����iP��~ue�j�fuN�]%v��Ъ-���<�����V����F��p§���:A���jG)����x`�� �7���X|����U$�x(o��{�@f�Bq�����ak�kI�3aE��,V��@�B��2��w*{��������4�:�.e��p�����~>=)o�$jx �5���K��*gP�K�.D���H��CR,'^2
�(7�"[�	2�}G�Us���KЃC�&�ݧ�Ga9���l���D��T��h�����	�=�')�<8��j�0���SO�2��-�DqL�7��0�K�F��-ѫ��D�cUS�O��X��f�h�ѳL&�U�a�f��ƺ���(��W%�a� B^9��/���8�����TrZx�QU��y9d�Q��hqO�x�z��j�mU��QSR�ۭ���B�|p2����u�<�B����w��R����x:�?䘾Ϫ���x�L8�0i�#l� �Q�B"%N�urr2l���^A�u��p������P��P?���I(#ɘ5CΟh�X�6�E0+<6��"W���P� ����d�Ҽ���?��P�vY���nȅ������#��;���>����=���^��M��8?n�?���o��[�e銹��g���0�miQ'}��_4�Z*��u!T�\T�.I��X)��D��q_w��8W����S�rA6M~��i���T���$�p�ic�Oa9i��{�UL�Q,;��x��ً��Q�d�f ��ꑓĺ~l�?���4i�/c,P��\-����f�������U$������U��&�-��S�)�%��yJ{����2�Ԭ��i0Rq�0ЫZ�6q9�FFzB�Ն9���\�o� �3]���)�9Q�^#U��%S�j,�JU@���'b��\ �`=6 ..n`����҉�6gS��x_t���ǵ�m�g %Jw��w�l�y掂���E�@6v0��3��0l�)���*߉!/�*��d�64�0�[U�Wr$1!u�0�*���!y�p�w���*,�*��|X�W�v�/��JR��t��D��i����tڜ~&d����ݷ6�jcy��{j?� c�D=��+Fs��䒷�&�+s������Ϳ0oV���������"�:��ƾot��4���X�j�.G�lU�u*�"��i�v���^�9���ž�kFLN�ž�NFX��2�mj�[�o;��l=�g���Y醇��_�,,%�_��>�mB��_�����BH����T-^���޻�=_�.���O^`k,/����v���k]D�LO�ڰ �={V9�a�0P��y�0s0z`��6?S>�=�Ë��Z J6$؞:�5ڷ���c�Z|���ňi�Z�r#���{��:�V�b�#�6�Dc�� KQ�[ncq�p�ަL���)���"��҉�LU
Y�-�	fM��:B��i��R"�@�~x0�GÙ���Y͡��ʘ�d���HFqz�U�ܑ3���k3��x<N%$([��b��  ���Ct{���ē�p��%g�|�LM>n�����f����\PJ(�v�P���3֦���r��G?k:���� 8�Q����s{oM�������Ҫ&me;��衝���'.Y��T4>Q��v��uٴ���y�4_�����q�on�"}��tvu��ۼ��{ ���<�"��`o��>!Q���45S �k}��I>s8�KV)�H%B�e���U'O���������05����xc�57�G��!���U!B��z<��F
2�D����^�[K�!�� �b�5�:�l|`�R�+$�RM��4MN%dҖ�f�c�U� ,�R��[��Ɠ�"
[7V���a3	RK�ՠ!��B�=5��s~�z�~��.i+D`�Q`��'Wq���kǷ��C�En�����Uzx*�.�%��v��*` 6~�*��6��Udb|���]Ȯ�1�e�������(���5� H���:�!I�k�{��B�wpD��K>�
l��D��{s0���#���y����m�Y�?�U���+������î�na �hU���/c������mc��Lm$*��K?g>M�Ç���d)X(I(���(��Ô14u�R��J^��]/Ğ�&�49P�ZxF�U���{Wl'��Ɵ��/W�l|�G�.��pC薜�N%`I�%��	53MUē���6��.�<i�=�*QV��[�v�hP��>�0���V���HKb�z����F�x�OI����hD`��A�� �P���n�*��t�����r=`�Sx:"c������lz�[֤/�I��)����`�,m������jL=�$\Q���{gS6$�k��?���,�$�[�(�8�cS��˕�	�D4��#�� ��[�R'C]xN�:SإCF��b���W壬��X���I끂�,~��׶�iy���D�Hdf|����$g����`c��#x2�4H�%mJ��&���;�7��H�����pN5�m���Er��9�(+XIdR}-BM�T/����q�h�G��@&��4����V����ΖVX_���3_���N�w�|�����|va�m�?�x���f���p�����7+�����΂���W��[HA�����ޘ���uf@R'
|��޲(��$�1�7��߾����N���9���<�0k8���<YXw�Bp�%;J�7̟�U�I#q87���c����tQ@vg�����|NMY�
z/��a���R�Ir/��i�s������y{5��	�-QRh�+���S�~i�;"�_�t0xm��T(�u�{j�kuB+2C�d����09�e����0�1�wo���q}g�I �ڱi�A��f�ݮܧ$��ct���{(�c��1��3�cc8��
��w�GC�`Ҫ���o���3lR�����M����wS6+0DH��kEO}���'��et.��"���%o8�Z참�p���Jl��}��|Y%M�ZQͫSh�G(bw�E���Q��hғ�K(�I�VQh����Hy��w��1��i�
=�+�@�L��C��C��.�ۯK�惛J�*��̇��#����{S!>��e�ʡ��	mt��1�.kD�>*|
���ϲ���5�>�y����)4�ƤQ�����&�l���-���@�3�f�h�C,�5R��Pl��C���'�v|��~�K�$R	�N�.�ɽǅ�쏬Ln�jP�X�I~�bn��M��S�K�����qnݢSk%����3+�Ւ!#[k������nm��ʋ�	N�������!m��� �6�M.a������
�T��8Oh�[o��kZ����>s�:|o��	ߕ�	�� �f����J3aX���ї'#�Pr�(�:f�=%����(Y#��䨯��vr#-[�����K��a)�pR����-1;f�fKN��kn+�7k. �%���G�r*�O��~@��S�����An����_�֦�x[e~��� �i�r�:�f�E���y ��E���OfS��	��bRJ�w'�:x �r����	�S�S5���cό�Y���,'���7]·�����w��w��*��/�*��Re���jD++�|��Ә��k��^�V �"���?,�op�Mtؠ�Q��~㮹T��;�%�.���@��sA�ݓ�F"��6���α;3P������͇y]޼}3�z���v�_�:Cl�c�_֎�����6Qӭv}2�	�2���+Zh'�#��f����k.�imO��_͍ػ\؉�ŁRU��¥�;$H�U2�{
8J����O$����	yci�������҈'=�y��ǟpe>��f�n<��vM�F�k����j�iCp28'���c�����Q�',�a�_��;2}�����<�uϿ��=`���;��3���[����C�q
i�O�Hw+�8.;�7��L�������<�ZRS �%��y��������2�3���?5G��HINݠ�t"K���X5��p�3=��uI�����{���_V� z\<��@�O05��	���iX>Vb�G�nȨ���H�0�[�c�J˸��Pl`��ߣ�"�օ:h��.��l@+�V�Y�͏�/1đ����v*+B�dK C��y�\3����/iU���8E&M
���DWI{�)@�Q�&�	"	�0EܞCQgB/�c���P���/+�>8.x,��X���%��!M5�/I�쳚�͔��fE@.h8�l�*B<��VG����0 ���Ǳ������0�7j�� e��Q��l'W�YF�J�><�����'$K!?���߫�_�Z�@��TKW:#�g����{,�Q���M�l)��c�n���AGo�!�x����h�Ct�Fψ����6� ~>�� 	N�*Q�1�U�8���sVD�� ���~�o��d_9rT�0}U� oM�[pY\����;	4��F�l<�[� �Ʈ��_;
70~�T�!i� *�?�i��ʸ:�h��iy��:8 �u~����Se=^Ii�����3�Acd���}��SGs�;*#ojX�D�[z6{�6��R�ˏtK�9s�G�qQ���y�����IS�i�PAĊY�@���i�PN�	�0t?Q���:��6-���a���4Sz�un�I$�9�u�Ke�N�I	�\����\�r�o�Ɍ9�͒v���W� ��n�CU]�V�tE���]���T��`������k/�V~Y���JA�갵"�u������+-��$����V0qh�`��2ie��&9��O��PJ����x;,�Z%s�4o
fm�H�h�[e�����= �p)w,����j@/^/SR�tU�Ժ|`J��N����ș�l�oI����LϚ�XY������o�"��d]��Ȯ�1�?�&Q���~�~����G6�oQ[�0P�gC�|ρ
��n����G������o����j_�X�-S6�H�1&2q,�w�P*�-O�EM��L�v�R"o���8�ZV��L�����@c��=G��V���[���1�"��n!�2�����3cA�ф����%��Y��l�	�M�;��{���=�L��ݭ .7r�CY��.贂DO�N�0�~�z�g-���CC�f�_���<�)P���t�N����X�N�zi S	�~��Hx�޶��E�qJ�q{�61�V�H�2q,hQ�x�4ķ�e���c9m�A��	K
�1>ƙ.[=@�w���E�\�s\7J$��4C<EL2�G.�d7\SKM��T8\�/o��˚w�SC��o�H
���x��F�k��$=]�f�#�����~�Z:Z\��	s+�o��XP��-���٠n^H/0� ��t(j�cs*��D���P�����C�wS�ْ����>�O[�u��+�mg��9Q@F�v�4]�C&!�ԽQ���cd���kq\:'|$�k;T/,]����'8�[w#G��T�?��?"��_B�a��,&3�TyZ��٦�a"tQϺW����`5�P�`�6v��4\�3`M��08j%.kC�lQA�V ������k�d��#�(`�'�'�W��eELymŕS
D^X�	K�V3�4�T~��5zx�l�u�>CY���`�*_~�@|pt�f�ׯv��K�d��VR�)�!����c.z��ޔk����d��a�ܽ��#c'�X��I��/�H��4��:�TN�&}4yMno���yܡ��A���M���<�a��5D��qw���[��-�'�pBp�{�����ي�$s�dܷ
��y��Q.ʫ���L⮆�Z��>7��+׷�����'�iЉ��W�3en	�����;Hȸ�c�Q������E4���_�1Po�W>��@�qI��w���3Rzzzj�-�1�K�K�3��e��u1 ��F]t�M*��GK������~�T/�֒�D��H􁟗�m	���z��R����\�CrmҤj�>ͤD����C���݇ �ꢘ�2X��O�F_H�W�` �=C��l��*��&{ҋ�?���R�(e�����O-��Zr���[�B���X~�s�N�.�gFL�Ҝ��v��	�Ն�X�	D�;�H�׼@�LĹ�L���ݨi�+��q�4�H;����w<[�{^	D����$|�L橨͙ �Vz�\��n�֥�=�8|�@}���RN� k���l.�cְ~��%�(F%���s�P.�&c2��-M��7-��aC��kǷv�2�[=Ћ���Y&h��m[ާ�����$��l홻��G5�h���+�_���o�R�'�t{9�RD	�.�[������g#d+�"Z�a��)z�̩R&=!Ƨ��{��ic��~!��2c�GX}� M%c���V���I�ϮnojB�Z�i2��`=.�$C��xWXO8IH�7'��K`�Ce�V��"ݶ����2�.����B�I�Ĭ%I���l�d��&�m2����E�z�w��O�Zl�
6�h0!{jgƎ��X�	���Rdy�a�6��'���Y\����A"�@;�c��a�(k�/�^[�_���l����
�w�C���i�ܳd�1s���S�$PO�Dg
/�Xf�&�5O��p7T
�@�Y�? _:�cL��M��E|l����]4\ W�^�7B]�d_95��{.]5��f9T�&~�'�H<�)��>�9�SWQ괓�֖��9e�4r�I	� ��	_����p_'���I��ka5����&�10T�~@/�V��% l�zH�::.G"je������|l���1���*C��Ǔ4E�N�$e[�������1�cJ�m�qCX A����jϬ0X}c���9z����]��z`����)�lp(�*�j; ��n��7�u�R�{���D+z�B���f�i�?_82Q��~�9в6����V�� 	���zc��A����n���/f�#?en�	#��
����oAzl���M�v�WU�nlt:2���Gx /%H�������=4?ߺ�?l}��q���)I_�hi�f;y���/���]H�IjaV�D$��W��&�x�vZ/
��eƔ~UXb#T uB0�YFF��\.�h�^�t�������~L�LrE��t��IR(�� )ĴGD��P7���
���>=7V�V�K�IUzd��ҁ`2|r7��I���7��{�տ>��ۆ(���{��7����%ʒ�`�.���ŀۃ���zej�p�nw����O.�}�`��/�}����.�p3mq���gm��&zBW�;����?�e��U�]_��y��B����f =�v�T�I ;3t�`����@�h�;ԋ��
t��������X����~�$����&�9���2b�Ⱦ(����}��M)�.pV����ނ��0*(�H���w&�D�}�O�+���}����졖kXq�RT�T*P��B��$� ��I+�R�C�z��ϥ>��'/��OrΑH���@Qk9�2KG��(T0���Є�½wmR�3���H�;-�xa&�ft_e"�R��]H��Ro]�Y�y笖7��~��i^�f�U3E{���Ϧ��-�cI��/�����LFj���ϹP����*��y�e<���[l���'����`iC��6�����L����6��÷����Fs��}�~l46�ƶ٨�m����ƶm۶�7ֳ���x���؝��s���#C+�k:�_0�.v�	��:��j<@w���GL22M���w>�]�R������ى���H���(X>���ɋ��EN;=����4�,�]Y��*MF��حLd�Q쫒���f���t��Uv"�q��l3�,�ngY�#9�1F��~�
��=C'��;���.8���wWbD9�,,;q���i�Ƨ�G;���/���љ��E���O��%�Dˑ�w'+��PR�Z&?v�d-AW|e�y�^����thn�ݜ��B���$�����$z����X|�f~�r��Cz�R�G�M�}��&F'_��7��ӹb׍��"���H�2z�V�@t�����/0{��ωV�R����$ŧ��^�<�t
��x�����r	x*p��y��ص]��_'��y��d���_�Ki��=�^z���:���r+��?��� �?{!V�M+��r�#'��L`��x�~JX;<��F�Ș�|��nX��!�@����`�q��E�HPrSf�n5��P��j{��  ��l�!A�r+����af6�͟�E�$�G�\T��v�Rl��\�m�גּ���PD��L�8�O�ڱ|��L2�}K3�lI�;�[f	,��C4��l��T����{ϓ-O���Y"0v�W`���OՆ�@sj��מ�����}^.��v�hB�&���J>��� Ԟ����\�w4����6&.m7ٰ��m���)��a �)�D�uo�q�Fa���s��w
	� �[�H�vGʍ~��B��<�~YS��������{�����)˾�(���o���̹�ܶI:�5��>_��W�L�W�4y�4(p�J2�!���e5yT�Y�hP�L��o��LzVA;�����Gd�ﶇι��Ʃ,��D�߲Z�VbB+~�kz1�����AAAA6�c,n >*X��c;!OXo]G;H����s�C��!@}�~��t��A�C�D����g�/#�v�ϒ)H<�d��K4<~'�ĨY�T���&���Wa+M��|K�:,V���	��^|��~�m��R�ݎ�b���{�f�N��cХu5??�����:;��$�*��R���C�F0�b#�vv���<=Q���7��ـ;��A��Eh��O&������כ������ �@�Y ��i�%Wɬ����ӣ��ˏSJ�PP��u~O��Q����o�@^_�+(p��L���� �(��=k���o��o����ө��7ݨ4�Kұ��M^>���+!G�����ɰ�5�#af���$Ƙ��&oBkW�z�K��89p`�l��U��~Q���۠�kMY4k��4�=�l~,�:E<׌�3Le�D��_�
�H
��SR�EN���s���n�I�,�e����V�>o*�a|�E:����4I��� 1WJ�`��I�v]b4hLc���Z��S"�p�����%�J��C`(_��	�<Ϝ_W����Ƥ���Z^P�l��hW��".��-�#�Az'o���tٔ��g�ԕ�-�`̸�a��ZX���Z�z��"�VCB�ޞ��m@5��]����i��o��ӯ��钦�ۯ�e +6D� )����z�/h��>P��?/�J��$ t><�'*��4����Sp�~x�1������~�������5�يk�N���w|�É�u7v�[�}\h���@"Ȁ�0��7O�A���}���I��n��-F�e��F�{}N�_:�ğ�-mK5V����&Ng6���e��2D+eC�*�*� Tiq��Y��e���� �fp��s��R��-f�W��<�˹��8�ӓ@��%���"G/�$+�5�p�\���-���1��lC=��)U!���IS'�F�!�hўP�o�Yn`y�&�$�ܒ�PUh�=F��T��P,�������_╩��Q"R�A��Q��E��ѳ����aK��=!��m�.���e�����������_ ��<"�,�"���]Z�3����ݧQ��$��d��`{mj�viD�d��}��H�i	G�ZO<,��ưQìg���k*� �ܹTF���w��c��W{-����"�T����赆[�'��l���bu�t��w
��|�R)ZzIb��F�C�٤"�:�77��ڡ�����P#:^_�27�����u�fr6��?�OT��3���]�a�`��k �����%��m�jv
���Q���yWװ*��üD]FQhi/��g�` �q�*��f\C(wP՜*sݽK����g�S��Ү�ƴa��	Rm8}���'�T���#/ݹ&�Z��^�y������p�,�n�n��T����o�����3�"�0��ۚ+)�GQ�/��>'�o'|u��-Iu䚻�>����Wu������0;��2�F�g�}�'�`&sxw�	y5w5��WE�i�:k#�{��Svb1G{h�Y@�a�#2���0��W��f[�>y��-�|�}fz����{��O���*3s���Z�yp؏�7�,_�������*j)��Xꊯ�]du� �B@@Q�a̾�U-�X�@v�s��`�}�;鵶�������L�sa7m��ų�	���ժj�j؝ivţta|jv�Q�S���E��:~p�����5u!���d�f���Tw�aY˼9�WO��ǒ�֛�Z�»�\ww֛�
�+٣���"56�M>$3W���Dr+�*��\�Zǭ8&�l�FVyL�[��a�A[���s�F��Pۃ�U���㔎��T�?e`x�Ń#���vN4���VB��R��Ԓ.Bgk9�xoR��������k��-���E.��l�*��Ӊ=�xz؂�]���W*	�������Ǟ�PT���j���C:�oқ�$5]��A�����)�҄ٞ<��/��r���_�S#�$�xT���gܯ��8�i�t�Y�'M����i���(�:��pU7���33���"�7k�.V��v��8��\��Q���vus�:�H�o"{?_�
��>t(Q>�SR\x���"L&��p��=���nmک;*��(?8��n62@�m�!����6�h�����8�Ll�%ҝOݍZα	ϺBƄ	�~mQCa���l��Kas>8F��L/-Ò3��}�X]n��Ҷ�����\�ŅW��>7����O��Z�8���%���]����xط469��]��.
�+���e��)X��I �Y�Ay�!���$��j�x�b�7G;%6���LZ���A� �(���z�j�<�00i�~�}�Y-���|�=L��Օg%�������=Ȟ�9D-�%�Ԅ�͂(Y�=�y�=��َ��	��۽[�o���ր��~�.o<�-��6u�N�ۥ��p�S��6�*Č�M�aU$�*�[�����7�sƑ'�~�};\�?d��q�S�E�EZ�N����������Ign�8��Ög�ϕ&o.��@W�5��y�d�jj���Ƶo4�K��w� �͔�J�N�x��_���/�r�nላC�"�6����$Ax�2Ɵ�$azk"?�joe䫘R���ۡ��s��6H8��jZ����9��$@"�!������
��lg,ꉟH�Y��k�Z�Iaŷw��Z�I��ǵmʲ�:ϸK����C�X�=�\�L�YJޭK��z�b��k�r��xib_u4�-��T*/\b��P���E/&�w,̰[uAq��N�赧���/��SU̨�е��?S�b��#/_M�
�;���f�=WML�ǟi�p:J�������,�c{"�#Kɒ.���S�[��)e��T�_єml��������i3����+�LT�:@)��s�q�9J���dg�X��߯k��)D`H�is��D����T/�^m�S?�sv�U�ᠻr?Bn]���2q��Z
��ҵ|��6$ցg�� Q���rh���~��˶L(i�{�t����UݰJ�2LO�[�&���lW�%3������2)r�*PW�ڜ��jp�y�ى��l-^�"�?�"��'��5��Qd�������V�p�N�4A<�zW|��{v�uu�&���G�Y�Ƚ�a�����51�9.go����z0"*�������.9�,]�:�^��ˤ���8n抠k�>�����
'=��'M���0�
��g����oH	�
��`�S5յV���䐳/��!�"�w`b����v)��z=���0�*	v����K;�<����Y�����P�eh@6gDT~l{�]���&J�g�;�[nś2zvP�����l%�����}A���J3-J\$y��b�y���RА
;t�]<x�5g�;��9t��OI.R�[d���nrՒ���B������-����.��X�N4i������39%L�n9�]�	)�{.�V����;z�h��*������m��9����R�7b�����>9�-~Z�/�P\jn������
����1ő�sD񗑻�!���>�݃F�/�X�*8���]��_��/3r�1gm��a<_�B���g���u�9�0�R~�W�d��������kD���K#u���;�*�
+����R���K̈�ͳi�����)�����!�O3b�����>N��H9�˭��`n�G�u���Pʡ�B��m ��5�Q�m�y�t����@�A*�8R=|�П���;��k2@��xZ��D�|g��ۜ�swצ�R�S:|��v�X���DJ]�o��:;k:�̚&�2��z+�Ҕ��"f(#�r*�TZ�l%���z�,����ֽn�#�I��z-K���{&j��q����h�){�H��vX\L���f�0�y�8_���j5������.��p7Z�����k���qh�v]�Z������}���-Y����c��.�}�Uӷ.�(�M���������A�����o�!�4�X[ҽ˱N�tY�(9}�k�%��D�wXݬx�����:e")���t>�:Dw�5P>1��o�f��R4�~� ���Ƴ��|	�|c�B9�zbe�@X@9A�{���z�y��G/����Q�ˁ��(LM�-��?�;�%�?�Jrmu5lP�mb��i)����RŁ���DWR5h������ >ZH��Xa\iv�y�/MX�h�b���<�"Az���{�Ŧ��}�3W����eA���,:|e�T�"
�g [��<�����l�L��w�;�ӛ؎S�MG�%���l�s�	�����cr0����V+c��㭶�8q��P9%��-���kWMX�P��W�D��?^�� ��E���n91~�@(x�-�獳�lRV�e��!���Lc��Ж�Tt���IY���������7΋5WI�Mf�w����t�y!�Y��Zhʜ**i_8��\gO��K���}9��3o�90Ρ�1ky����ph<J�'pF|X�cM� N���Ϣ-���z���X[ɥ��
i�N����M�g�!��6S���O�0��M3>B��Z�:�+9@�c�Kh���6{L�j8O|��#��J�u�:��b�Z4�(����0��^���pU��]��+��J���k&�[Ĕ�	QT��X.9R�r�lfkMH�yB�
s�H>������ڜ�Ewr��J�EcPc������7�`��Iv�� �)-���UۣL��G�d�)U�ּr�ʋ�	U7�t��*zo���Q'Yﯟ��{86-?�1B���%>>�㹳M��)�(���+K�GQ�d�8HԬjO<lX]q�]Fr�~�D����:�؇2�����y丛��w����s3��w��ƙm����7�~C�|aA�UgǛ�!M%�N����B0�ֻU7`��cR{��
�ca��\1]x��rش��B�ʴĖ{ӥB�ҪƔlج`c�\4�ū�-��a���l�YBU���L�u��ܸx�O�|8������&���Z4Z�l9Cw��J���Z$إ@i�63,}?�vY�op0A���0nۂ��Ǣ�THW����@*����Xv4?H�+]�^W �B8?ꡮ�.�݅�`mv��m��=��X�?6k1�s���K��b�y�qb�Ol�l8>�<�S���_Rw"&�7����AIX2�
��qv�;��:R��Zv�w�񽌨Tz��s7Z��!a��.��p���W�O��7���5]~���&MIs|���x8���'�}ju�5��qDA�&PW������Z�=�B��Bϳ������i� ��I/��x5	nH���4���[.VR	�ڏ�}�X��m��FK��|B��όf������@C�m�x��{<�1ə*���-�s�䯄�qSڗ�\�d�N���ߗq1Q��F�D�����&wF�S �D��X��������׭�#UڐyK�����jBK-��}���Zx�z�z�f�K�B	�ޞ�ȏ��\�������e�M�3"�' !"��2L<e2�P<�ƛױ=�>�R�2)4��ފ��+��0���N����B��>1������}�"G��͸Y�qQ^@��PN1(j��F^^�eDI湶(����gI.��11����7�Ք�@SEU}vf��]��$�)�l�4��2�3]�M@պi�R�6�Pc^w�4�r-���^�VA	sጝ2���#U}��zf٥�<.V�Gw0g�M^*Ķ[LI�5 �^�Y [U}z�_/j��D���)Z}��m��k�u�KPw�lv�l	^FL|�8�c~}[�޲ƅ7��bW4�B!!m�+懨�_�J�h.��\S��3Cn��,�ɗט>��x~���|��z�	=���v��R��DY��4 �����	��;��M����[�5�QE��4M�=hj��>KР�#���\����TaU�D~߻�1B��I��Zd�N2Ї��|����Syij,�Wvߗϧ~��(�0>�yg��8yV&5<"���Y�裠|�T�f����@e�'��ݮ�ڞGءU� � ��W�-(�ؑ�;�х�y悟-�qg.x	"�S�i5�W��A�3f�B�z �~����k��]�u�te�fa\bk*E�#���>X������óY"���ġAFl��Aűج�&0\�揺��hK���c'`��U3.��}٢�){cC'l30��L���J�����&'J>uS3M��U��y��f��u�$�ue��I��t�tNl�U�;��_ʑF\�� \�P�y ��������v_z%V�m>��j���x������@�v�`E3��?�^<Hf�������Z��.[]��
�����ْ�F�2S,T�~?��]��ŭ't
�a��aQ�	÷v���+���>1и3B��dK��-�����+qw�]σ�r�6�^Aåo���8M���|;�@�~���+�Mr@�{h��:�~�@�h����IIz�_�!�L���P8U���fȮ���A�WZ�Q&�7��1�a�%��i��%o�PEK1a[b}�sּ��h{�VD��Z3��MN�� ����%�o�5Qz��/��Lr)�^ͼ��o&��7��B���T[��1��@�U?�=R��y��
d����ɚ>dɞR��U�z��:����-�}���HX��y'��I(��is�,���o���>n�P�Ȯ}����'��oe�)A����<f!�0�3D޼e�g��b�a��Zn�+�%�r��� ����xAO��������ՙ��� F�����WdG�NNcŅ�7���8���F{���*J��#T�n�"V�Ӗ� �H������ݳ����pi�NA���G����X��[aAH(m�mcnU|jS��S\y�怫7��_I.����nn�r������.��I�#���E�Ųap��~7$��ly���{�F`d ��N�D�d��rk���8_VY��~ĐK���2�oZ��D�y���J���#�����p����0�ɑ�=E����2��9���D�ؔ���N���Ġ���'9B�V��k����HYݤf�bi�p�]����c��~�^(,G8mV�鳌�� g���J} b�,�bվ;r6�3�ӂ�K�M�]Դ�-Ԝz���R�Dܡ����Y�i�ȥy�D� 4�����+[�tf�q;�l���M�U�	K��\�ԑ��uȍ��d�����.iA)��e�1 g<��*I.�4MF��}?�*�=A#�(�=���,��@V��9 �g� �8��9φ8�p*@�,
j�O��?�
6y���c��8\1�}�gx���r�_��,�5v�An{��d姧R�Z樅%i跤��BW�[`Z)2=��r��;���U�_�/��\�g&��Ut����+
��Xv�����i���4���V5�޻��������9�qQ����]��{Ľ[����ND��EB=�|���ZM��Ж��:c%^6i��O.��0C�����!����K��~��eE�w;l��t}�L���͍U�B_�) /�
[���OUP�n���Q�)�L���(�����V���>�d���پ�9|��M�����{�R��Oy�x�(}.9�����u��3U����7���#��z2`K�،2�D��1�W��1�)��x\#w��AE��xo�����YSG��T���"�`�0�c>G�u[�hhDh��Pʹq��*��
�<��<�H�w�f48��L�h�@cW���&{�kI�����bC(�t�&'=SZ�\r�MZ����XPgt�gZb���`r��3L����Q�=�4㋒/��}ߋ�V��S����앶�<�(T�T�*�kHO�Eԏ�~@���{O�2W�����%b�v���KP�~X������?Pz���-l�G�wY����c�C�>#��1��O����f!+�����~�&{�����Y]�q�v"%yY\��X ��2W�]�IotH�������;-�c��j�$�>�� �l�z�I�X�b]�l��v���j�pR{�#(! ,���3�;졛yz�Rn���vL��c��u�����֋o:;�(R�L@sQB^�.G-�����s�����t����� ��)���s^@Cx������WWo��d��<O�����(���������E�_.,$�D�����un��E��k�����X󓘀�)Sm�����t|+q�y��E����G���-���wD�� ���ۄ�����������n��b8}�3�]�x����vrm������7o�����65l?E���!d[���8���+By@}]W\e�{�z�����g��?���/���~"V�_���5�:�h�5�$@R�D�f,�O{ʂ���6��,���,3S�����)<Ob�׽!y��f&|3\�EX�R7�$��آ-�gw��vE͖���.���Uu�M��lr����ۿf,�k�V�Q����-���D�� �ej���eSLӂ2�	�����c�����x֔�Y��[7����8��߲ !�G�"'쵂��WC�'�ǥ���vΚ�oMk�ġL�5�J��H�b�l�9��q�Q��!�eWF��啎l=�e$3�1/bb���Do	�/�ٰ�Vo����/~���m��rW�����C��6kz�����D�e瀳�g^GT�-H��/��,�����3̗ڪ���5��m��L�_�g�����͘U��M���`^�U�	9D�>nY���~�+`���T��y���x�T���Z��44���0�ut�R�\P��B rHSa��q�!�H�D$�*G���־}#��5���o�0���h�^����RRE�2_^�:���ߣM���u	2,�)���=�s�s*K��A�9,�<>���8��1L��+?��'�s�*�J�'d��Tq�����\hgQ��lK��RZ�����Y����� v�`ђzft��3{	�mEf_�ԡ|�����9��ʘ8��#���'�c����
�S�aoQ���Mf
ۥ�1�[�9RGT�~W+Q��:_��H(�Υr�G�AC�r��������	����>ȨV��Х�����WmX����A�f�#j����Isr�"]b�"v��7 +��f豋{��I�û�%�`����)���e4,�<,�SG&sV����0v�/�;���
�9����9�3:��g�������[+�)���3�%���;�3�^�7��{18sl��? o.����pЅ�r=��M?���R-,n�~�z![6y�i�o7�U�)��c�D.mg��ΐ��o���٪	��@�mv&�$ˬ�[��%QƖㅕ�F�v�BS��N�	7����u��2j����?7��-!r���9۟�Vxc%�on3�#e��f��&�`5��?�UەWu���6�2Ԗ�]�n�Z�[�����*a�����JI?>��E��r�3��ݸk�r[˒�B���5�3���9�U�2载�g���jt�d�􎋙�G��&`,��$jt�rr{�շ��>ᕢ]X!�����U�~����z�l���S�1X⪀�bE@�:|�i�uS>ǖ�V5+;�TB��GM�We;�.�ǮA�;{�K��=	����C������Yi1<`� �~�G�_���^L��xu0��g��)�K ��ՉKe��R�o�(�u�u�+���.ȓ#\���	#
4���@��T���S�iy�D�q*%�-���&����ɫ�lE;���9��Ǭ���N�k˓�������5�|Kc����U'���;Ϫo�7qR~����4�o����2=	l+�f�Pr?��~�Lfk��6ʬ�]�g��%�u�A��/��~K����=�ى��}G�z��?���2#?lw� f�nG=�4�7�+"��)q^����Lp�'z�U�������u��*��S�N�ބ4�M�(����V��^^�Ƞ���%�ZO*cw�d���"5Mh���-��W�m"�����$e���e����}`�f��[�,��o�y���=6�_^����ŭ:C��W��ջ���C�X�n��������m�,W����U�0z��a�gY!�"��.^T���{�^_����Dv��f�p�a�2��X��C�������ɾx�AŔ6tYYY�B�trx�z��Q�]d� G�Lv�"p�T��q��eo-��l�⮇��%vt��y	n���l���5o�%�Gt7����������r�������P�C���#���y�	̤'[-E r��҃fu.���ڭ��X�Opn;�j��ҕ!S�������1y}i�9�1�3c4|���ڪ�N&%���mu�>>�,Lb�0�Ti$Й7[e#����x�t���jo���/ꓷ%Y����Qd�Fkj��^���{���*v���뫣�n;Gu����i��q�;��
�2��דҧ�4��Uٔ�a�gL���l�lbJ}Ks�n���hG�Q}���yb��nf�v��֒g"W��<zƛ?�!�^؎�YI�l�~���\�dOc�ؼJ|.4;̈́e�ˋ����m���Y�
�΃��e0X=
���LG�] �oi���̬��;]�:4m���h�pQ���ǒOJ��I.>��}�P����R���[��`8R�*��{fYӵ[�t�4�k�ev�l���S�fCѵi���F����Իڧ���A~5/O�#��ڄ/�K��=��\�v	S�Ι��D5?� ���wm�N���;�W�vL�Z�g�����AlE�G�M��ң��D]�n�hx6�Y�� 	��=U4�2 �G"�Q V��F����#��!�!>��$�ԏ6!/O���.w�����ݶ0���W��o\w���ۋ�E/꾨���+�:2�D��4IԧF�#��A��&�}�;(�J�A�T7ۙ�'�W]�*9O���aL�~�Q�>�2�6ɵ�7g{��PV��l0�=���z���r�~��_I6�-��{�i�+ժT$U�P����za��{�V(���5�b#ޮ���i��@�k-���[��fňQ|��@���$�'"���`��Nǂ��5o�˜�,/й�^��K�߆	o�ݎf W�rj��O���&˔@�~0DI�D�֔�����)�)!�hc��ݵ"�wK-=u��(�ǎF�*�v��"���٬�#����ҙ�J�o�Q�BK�������3�:�ܪ����}b6/�"��Z(����N��	sZZ��9��웖Q�v��mb�\y�#c�T��;�A�~�!S�8ό3j���ļ���&�<4(��iV�O,��p��u�嶼�vS���g��k�T��.&::�c+� R�-�{��޽� �����tLx�`9b�v�$��L]D0��:��]A-�B��@�
�A^��0@������VK�tqߑ�r�����̈�aS��]qmh5�	��J��$�14�e�y,�SSZi�/u붚�+	s�g�Y�o;��c�M���	��󩌠	*W�LW��.�<P��-�aE����t�}��������w��8�Y���E��ˊQ7�a�?�IF,k<�������=^���8�p�+eb7ze=;���2��Y�&�%�;[b_��V�^fD�}h0s�v"gG�߈V��(N__��������B��FR(��:^:�>E��|��rP� �zJǅ���޾u�R�:� 8O��j�?�å	�>%�O��f+Z�L�GsT7����U�C�/�4 �X�!��jn~A׮Z�g��XjA�@��7��T�����R��i��J���в�e�����)=GJ���~SV��ui	���������JH���Kw�R������凉�z��L4}���B&hqf��k��g����6���2E����Y�)c?��W�z��MH����2�`G!���H�鹰�Y����%�-�4nkq5p�J�"-_�}#��h.��I�t�$:�1��v�����K��EI���A[X� �����}��57�%��mqE #@��VX�)F��T�y���5�D?���<��rNi�:��ޘ�\z������)xX���nغC������v.�E}>Ɨ�J�>>�W�tj	�N���V�MT%� ]�އ��l˟����H�iI�}��-��&ܯI���V�-|���ҕ��v�ÄH����X���\_�h2�0�~5(3Pf`847F3���l��y������	$�Uts����3S�ۂx�=?��@�s@tN�A��ѿ�we�~��k�z�^�h��W�2��.�23N�X)0T���r���}�X�Ȣ;n���j1h�b^ߗς��i�/j`�{i���Lr@�jh8�_ f'E�/%0����zJѣ�*� �,̸O��	�ϖ�fr����z���s�=���my��C����γ8�.G����a��FW6�v�Y�o��hVV5F�B����!�%���o������>�X��*|ڶ��e] � B>��:�z:YVL!��5+��5o�3��_{1�X8 �5�泀�;�TA�=���3�]��Ħ�|S�p�W�P�%]Z�am���AIS[Uy{j��h&�a|�hzx�A�<.T�:�cD���e��~�'�o i�mA�/�R���F_�~(�1̏�S��1L���葪��e��p�x*�P@k،cz�$����xy@"��8��o��v���I��+G����;d�ni.���a/�����fU����|�����xT#�,��E���/�+�=�G���!3��v��ьP�f&(�L=�^Um�Rή�F��e��M3;~���f�r�_
& �9�$1���KA��9���]r\\j���������HW�-̰�3[�i�Z�-�TT����H��푟9��Zh�,��)7ϰ���Մ�7���w/�^o�N��*�{�2�þ\�����_��hr�=Tr�8Z?��4����	p�޺*�ӝs�)e �Ŗu�+A�JI�|d�)o���1��A�2��p���+�)�����:M��ܺ՘�����~�;��
u\�~�f�f��T��/��[��B���m���ݝI�M�E�U$>{�	�#���>{εA�B�!����v# H�籴(v�)g�� �~��z� ��)���~^' ��,
���%x��d"y�L刃?B��QW'�A}�d+	�6!�x��'��4�|����1k����P�EA��)���{�t�	JB�:�6zK��#�O�2(�D�I"O�3�V���pv�J`N�nT�<���i*�Ul7�������'�6��L�R�����>n�1F�i=	����dR8�juz�ɶ̚%⃄j��MK�.h%�,SRH�0�^~,C�2���ō�v�윎D�_)���a�~���7c�G�ſ0n)�������p�(ޕKh�׋Rz�}]�6�4WV�rb�
aH�e�{��F$Iq{�U���2�oԑ�{�a�գח4�R�q���R��0��_�����CsJ�S�k��h�5,=��������Y��߯����h4�����������X��cz��8VŊ�*���o��$[�Lm������jMl��L���߭����w~}TE�9�5�h ��1�MS��Y��DY?C<�`�끔~�ݠ�̎@8��<�8|5fg˒923R˺A��<]��=��9Mw����>�������V��y�H�7�3o��mH� 9�ۓ��EU�� ������OU�݁��i��G��#d�8��Js�"����+U^�V"{v�������c-Ŗ�}��=�%A��9r�I��=:�x��߲Q�F���8��mgL�"����$��i�5���Ϥ����M>����'Qʗ[�f�)N��M������i�P��!����ac<��Δ���氧^˶�0ItΜ;NY)��P�g�0���R1'u�y�'V]�v�4��v�}�k�܀�5��Q9�����Y�,^��uv��hW1f��I�}vʗ��je�a#;��3��iרi.<FV���ꀵ��X �s>��n�S�qƂ?J����i��Kb���u�1I����MMˈ��p[�`��s|���蒭�����bK��V�J�~�8�������!R�;���u��X�T��A�F����A\b��iF��'����#�VI��7PA$�¥���yn�
K��#��"�ÉƱ�z\���"�7�h��1�E��侠��8�S	���"�'*�٧�BX�4%~pf���ו�Cvuz�{Cz�ɩ@H7_�{.%%2㸏z�6�2�w
$��՘\�����ڄ��-�yy��{��v^%
@`��2CP���d1p_��cP�%^��`nԞ�<r�*�aeVO�U���)?|�ܼO��o9b���_@�P�)F����A�nrD,�}��䫦�ma0$�W��8K�Z0�C��k�u�	��fJ�`�=�J!v%F��X[ɢ��-wd�!3��t�	3�s�=�T<$�Z���x?�K5�4q��9Dh8j#���0P�J�����´x�Ʈ��1���J��H'�W5�8�z~��>��|�aZخ�s�p4�R�R�:�$��ؙj$���?U{ms(�[[���=U�����[���Ә#�a�+��J:���_�j�A��y�=�r-j�v���y��o��������p̴
zO���4��E3#F#�n�4�j<@Z"G(�v*��ecLo�@Q����fȬ]��œA�.+_T��]�ͧ��~b���`�s���F:Mf��q���nQ�;~� G�C�x�t�gp��W�,g:��厈
����m���ړ/�Y\W�F�ﹴ�^(��k��7S�e�]�X0��@L�-oX���+��M.�[~B��Hdو�2�,�9����f�/6%�};�©�U0� _���V���BshП[�]3χ�6Ǯ��5f�`��%�k�����PH��0or��m�W��L�G��	��@�ߩ���s܊�`�_�V�;��f�m�L�2ΦkL��$O�J?�0`_��7�ѹK�"�"
�t*i�Ҧ���j��,.Sn��	��˺}mz:/��LC��W���F�8V�Ѳf�qI�ގi��Ф��ܴ��$a.@@�����u�pE��lA��k����M��V˷N�^�y:�߶����?��Jn$��X.5�E�5�F�����(�p���|=��@Ab��t��?r��Ш��A��,�hو�T�/�D���!��lص�
P�Iө	~��p��\7��\�MD��'��i|���iJ�~C=@-A�]�&	(V.w�9�h��f�ɗ���d�	��ٵ�P�����ݝp�K/�H5�o��0'����Xs`�I& �AI�ƍ�{.Rġ�ֵ`��S�t���9��c�rgK�|ߪ�����Ԡh㩬������(I|�Z۱ȁ��*���Ͽ�mN���)�vk�+�������
M��@r��7%̈9G!Q߰?E.�ٓ�;�d����}+�֖D%�FM��uLD�ѻA�2Z�:Z� j��>��DQFgD�3J0C�;��������{��s�Z����{��>�4�� �A��Np����>�g�!#��C�?��tSI`���m�58"Bkk��I�ed� �i~!����	<��0��������-K�洒��S&��q��4�'q�B��б��;��'�����6����S,ICam�N��W�o<�4g����s���QH���85�4Hn��W�M�?7ZB����j��:-C��^�,0�=�hI�xy��)S��"�|-���0Y�Y��	?m�#�_��ܮIr.�����p����m%�+��0�e1�$�WH�����>�,Y�|�0u�泄ӑpV�㓓��;m��k��x"w�\m�E�8
�Z�@Lk��^S.@�{��+�Ҏ�0��j��m�	����@�>�
�E[Ҙ�Y��2jx�gfqpG���"4�c�7�Ȩ1��o��)�uVu�m��a��CO�o��f��݃����6��Ӓ)��߀�J~��'�TBI})�%ua׏UW��/j�wK����y�$�e�95�/�G���I>���_s4nX:�k<��ݐf��zѝm��:���[�V�����ߨaM�Th��VtԞk�QV�Ό ��4��7���ju����Z��Љ�"�H�̮�O���N��Vɬ����[�> u�cp�v��~��֛��ک��{����ә�l�2"9���5[��V����Xy���zF���p�TZb�D3�r�[�߲�����Kl���W
�C��v5�� ƾ�Es~��.�|�{o��ҋ��Ƀ+����c���^��Tz`����[Yq,��x'o�!Jl�xL�{���*�Mubeuj-�_�f�k�������SD)���.���>p��BFm�z"�����Q���	U�[jf7Hgu��(�BS��L�y��lާ9��c�uks=x���$v��s�,��*|
����br����$|I�������"���a-���t"z�Gȁ�����{~c�����C��w��`a ��m���J�v��K_�K�/|���DN�����+=g�i3 �X{MTZ�F��m�K��YE���s���f�n4�I(�y�)�x�wڪ��f�M3$�ōP2<�oQ#O���DrA*�4 d�z�ց[)>
�V�2@6��q��o�9U���_}�&�
X��| kِ'T�h�RG���|��R�㸹|q�8[tGf��mǰU������5��o�g|6���5鴑j���V�g|�Z!�̷�Ƌoۆ��?źQȘ��ħ�5������V�}��:��m|4�v>H�?8���=��핃%��?u�S(�����o�%N�����S���������ͫ��%0��a�~��R�����^���;���VNK�{�xun��w�)�_���k�uh�� �r�^<�)~�g��&��<�(?'��?�����@����S�	�X��ϼ���f��l~``���<���C��Y�{"���a�膯�p��]��1�9�{^F����_�鯯k�X._�����J�jD��>��
�L�+�"U훾Xzm�J��?�H;Az�����5��cA(A]yla�x��\[�v;���yF��ϯ����s�/)؊��;4L��Xw�|<�-_[���x"zЎ~&8����"z��F�����!	#W*����5D�	�&� �FEX-d�ٯq������f"���{SU�F�PWw�]��dM
���r�S^���w�Y�����߇�4Zih�3e�Y��1�
໅��?J���\8�-���%f,JSI�X5'�hf��~?����	e�[)[�z���q�Nl�ȧ�8�J!��$�R�>��\�������u��!]�ֈ2��Gv�ӃoBd�QD>	G�aց�~ p�c�D������L�!e�l�6�{���T}�q7�L�_퓚��X��&�;7��G���#@��	k�_I{V��ˡ���$��I��2u߁֮��{��qu)�U鳕�s�|�Dr���{/l5�����k#z ��v;hn��xļxP��Jͼ(���|
����/�)��w���`�G
?��pǂ6����jB��;ў�&}�kj���G�ʤ$-Ăj�(B�M�L��~rz1��(K��{}T�u��m����>{�a�\a���W�S3�cl����$�N8�7����b�������Wţ����8�N�nE�i�;��)�G���$D���aK��P����w��.U���}�㤡�q�x5.H��)u���p?u�"�����x����n���a�ۚ����*7B�I�?9�~�V\��9���8"�/@���}�޸*~��6v5�_d����1M�tOor��%�1Z���T�l ��s r���Rɳ�[��O?xs���7;�l���s��&��?�Pa:������'_9g���QK��
��-o堤g���������k L�R����t�����> "�������"k6\�M磧f��ޮ���ƯW��X�)�.w�+���V����������;p��ji����)��zu����p�&u�D��b���ҹΊ�Zk�==�n+ޕU+ 2�{vd7t�e*�4�'����رF./�C��7�&�:Q��9�zTl$]���F������.�HLJl�b|n'�lk�wyOT��޷�8��b,u�W_eBZ]?�Re`��˦~����;�Tw=��z ����F�h#n.�����獪<�\�ď���]
!T�#4Jo*b���նC�_ޓ�MS�o�&�p޸��!�w0�"W#?jy(��E2�3��Ņ�4*J�>�a�?�|@FA�T"*���f�
h���eL(���<"��6nb�oH�~���#z��N���'.t�gGx��T1Mi���D}�θ��KD6�4�(�mo��?���䍤��/!o���]���=�D�7��
�9(���Ц��Ajq�ԁDY�^E�|�\��.;��\�$;�5���Dt��͸CS��0 >i?�}~�kϙꢐ��.�b�qj�����m�������ޛRCr�İ�i8OV�H��w���b����6���-�*;�
�G� ��on�@�+Ǘ���@k�¶# M��\��[�(<gb�s�4L�NgQ�?���f�eP��۶��=&������j���C"���~5�Z�ݥ�{��!��G�@(''wKI��>��3���� ��їg������.B�7��O�kڼMj�M��G u�b��(vv��iz�+�E�I�ʐ�U�n���N�
���������h�n1�n0�A�	��nᔱ�#���\�߅�����d�y����^茲sfh�\���������H�ۋ�M���Χ�g1��(K�3gF#m�?�}#/���kʛL��~��Γ����9!jh{Nf��@�:�1/��[�̽&[���'8���s���O����s4�(c�.�!�fX�s�W�`�R*�F,x:�+�z]+�(�-��>����Ǻ���"��9��_*���6D�0��^:S���(s�s;>R��(�H�7��X��N0hґpa;��Yu���$������K�}בO��!�����2�u	Q��i�}S��mM�ˍ�Y|���~{?��o��v�ˏ�'�Gv:vT���{K��N��Ǻ��x�}���'��Υ%������I��5�;�!���j�O��+�O���ZY����V$]�>�ƒ�G!:��m�eR�#��1������B%��j�c^����*Cj�n^���O���5���)n��T��ر�^��,��cr����ص�b[�\vz�/va2��~��a����������K���Ug�kٔx�{� �&�e�˞辜_2i�������N�l�Xc΀<�%1�<,z޴���A�'����,��=ؖ)%��3(+6�+4h��HƑl�誒�?�E�c#�]ݶ���Y�Q&a�C�F,}�x:P���X^�>~��Z���Gq��e��w�{/P��0�ùJ辎���}�X����S�����%"�h���5(�!���c`�ʬ<��	���}�F�����@m��!wx�#9�n��K����˙�Z�'�u��uY��ɦe �o�1.�e�uLys�Q���g�}r#6-�"�O'(�����fר/���V�x@���u��q�Ԓf2��S�y����Ѱ�X�W\� �c+�V�1��s⭞q	|5o%��qJ�6/���:��p���џ��y��u�'RK�z��*<)���V��L٠9>aAµ��T�^�
�7PG�;�����va7�ɖ��ߚ۪���@%�t�>.p�>S^��������Ⱥ���2x�딬��j�~����2����4U�qı�����7�hD�N�
p�%\��]�A�X��(���c���}v��E�^��Bt�(��l jG�펭���n���N)�s��wXn�ܰ^���mn�v�)1��c����՛��{�W%y�{�c�b _ ���8X����V�G�]>˷c�x	�����+�y���K8���ik裿��'���?�R5�)�~�]���"����:��x�
Ұ��U�u��c
�
Fm{Lma�̟g��;�n����Ɩ/��!�W�!����0Y�2��!;-����4��Yw�a謀��SQ_��e��Rǎ�̴�����p�+�|Q�B"�0�r:�n�<�A��N䭾���:�-%j���"b4�� �/�X�P��SSy�t𼄤���5�9��C�Y� W[@X���-�)�h|	��Eʨ��$:�G9Ywdm��� ��I��B�]�M
�wP��$0�V���L:Ê�K6�mы�7���QK��
�J)5e�h�-,�%*5�;UE� �g����*(X�z�5��߈�Jq8��1F%i����G��%�n��?��h�1�����!8�h�d5*o��_94B�d_j���V�;$����>�<�`Q��-K�c�>M��6Z	S��g)ʡ|H"}����2&��.�}��z?lM4���h[�s�/IV(����'j��O����߭��#�����`��bi�7,QK�{ޞ3�������[IA�4S��N��ib�v���v�ʳڶ#\43�o�!��ދ���`H�����}lnZC�]��:+��Dԑ�\�239⸆��v�tӋ�fAy;�6��=�l��-Z�hlz�/��lS�v�,���O�9����v,s�����8��L�
��b��@ۚ��|�)��g|�z����{�����BU�9����U��͵�'@\��m%e���IC8�~�nE��;8��	;[;�`qW���)���c���9!f��?
��㽊U,T��Dj�hFX�?7����b]Ǖ���b��W����x��~��͎|xM��p��>���e|&�٬�T}�*�����2����LX(�r%�:7�eYC�e���&^BU�����=�Ss��W;F�6�:|4k
isuL����[�I�b=��*��RM�y�rw�'��,����(4l�����ڞiQ; w���$��FH�;�b(����#��K���R6;pT̈́Uwp�H�`׀z-�N���z#>syr�46 ��jq�l�L"W��Oojə^=�ګeGK� ;�2ܮ��JX�GonU�G5ӊV!���u��+���PAV��8)ɤ�s��_\S�q=��XwC���e�ږ�7||j`}	�L���$�U�h#M�aP��3����~�继㵂'���_�揦kN�mu�.�Z��V�e�~%4<P�w{���E(���c���b�yo,+4�ُ(ΘxXJ;(������d��V�����nP�L���BL���\�3��FN�,ǱY�"�M��}{�Fy!�����c�c`�X�z0��f6�|��ri��/���_��&rPѥ]Lw|�2�]�����d���	������Xm#b�\��T����N�mlüO2XW�ZVʿT
�1&j�� ����,p��M�L�V�ގ':v�$��Z����e~6t�Eu�P$S��Ɋr��� }�tr�e�U5
�K�W�5�$KԪ����E�V�`��k-J?���;�o�M7�g���c��8�IT��ŝ�����1	^���T������}���қ��* �/�a2Y�[���i���&�2��o���k�j����������f���^)�v���B�|l�C&j�\���Ng�1I>��>�r��+6 
mg����njp�	:x��A��P�eK��吕����
�Pd��֡`�j��O��n��鎾l��z��!�M�Ck�'*��y��}���ܼ,5B�����m�_|9ife.�kM�y?���x*��}{���N�t��ѤWy�zC�c}� �i׽:�ic��T��G#|I	�|�zP^B�0�9B���F�;�b�Ւ���g�.�x��j�3/8lOj�u7���-^E�r<&z3b�!cY�3�c��rǐٮ��k/ѥtl�~~���:����O`c>Ϩ_��	�s�~^�0W��K�A�wò�,j�$��jd4@��<:�V���V��e��^xQ�\�>lF��g��Ur 
a1]�/9�.�4vB M '.~�8�8Um�т����f�ZL��*> �~����PY�&��y�r?���Jm=� ֲ�M�lO�̪���1��x�y��ǟ���M�D�	��|E�S����n	I�U�wIАP���5�6	�3C�_�yw�a�Y3���ʟ�c�
��*[�,��@���yu3���_������,/�-%Ou`�(Qez��5�!Z}ʹ�,�V0 ,8��܁x��^�ȹ+Ӓ��|}��Z�4jD��ĦP���hQ+�n<o߸@c�o����.M����'����Y9�Ϝ���Xs�$��Z�H�p9�n��������t���~�y�)q�ѱ.��ͱg��nZQ�1����d��v3�������`�.�f�'A�W>�\��\ts+В[��__%O�"�WV��4�62��5l>\�P��š\s+$w��3,��E�����AT�S�΃�i�P��6�Uzmf�_,8�bI��C�h�����>CY�;�*䘲���	�%�N�W�1��\�ҋ[t?�n�7YX�	܉o�΀w�����5gv'N�޻kJ�T�%�(�p�tę"��Hj:z�nGs��4qJ�W���!<�1Ŗ�����&�r�~R�bI�ت/.���-C��5���6�2����p���bDΰ��)�(�X��,B��c_gfH��<,���\���lw�"���ӳơH�Й��f�c��;B�懅���� ���<�bY��?[�K.A�պL^�U��Ap��D� �i�D�Nc����� �fu[�z>:傀��*�GHD�D3�Lmq�+����tU&�YH3Bb��X�4uu��Tߗ4���y���&��)�V��M镋�;,M���$�������s�i�tǈݶ�j)E1f�t��.p�N��m23a���.5�:�/�%f+���;a_�Ș�4�q0�n�lu|N��}��hOL��}Q��x��V����M�d�zv@,�lKEy�<[K���,�f�u=�$���x��9�Ւ^�g 2�=�>�E�j��
���$:��(Rp K�x�v�l��[Ph��s�R��T��_��W��ø�n�1�!1I@X�w�@�o^t�yZ}�tdb_���$n����`�$..K��M�é�/�*��]
!'���:�\�Hм�xL�-�
X�����9���ڐY�t���`P_\���r��,��vJ|%]K4�s���q'l��������჻t��DT��g9�6�rp򉿚5���ne��طpX�|����O����녩W*(��؍;�u�?��f�����#5��и��b��6�.�C3]ݖ���?|p��%~��>�_���.$�����*�s�?����l��I�!��(��2}����d������|b��hR�:�ů��{��X
n��7�#Y&X<�))=X� I��$b�Oej��f/L�2��5c�ot��L�b��{#(<����ӗ�y�����<.�<��j��|+4o9�򋬻���l<�¯�u#�p"�z��csʆ�,Y2���B��[���uP��r�x���"|�4��H�b��ƃ"ڹ����KG���36ԋU'����me�]��q.X����)�^%{z��r22���*�T�fǢps�S~�U�Ž�D x*��O1�b[�ς2z|�|��&�.=�!v�p����`м�c�X��j᷷��Ϟ*�9�ܪ�
�r���\{@��.�eQ:��17/	�(o���g�m�<�W���L�y����VMقfPKT���;��.)OϿ�!�����[����"�����L��+�������޿OɞF��u�j����3�*d��Y�S���������222��G�F��&�"�U{�����(?̅����������7[��O?����/uۻ���t����VB�)|�!A:�{�W�����[�$��j�0y�J�/Us��)͙�PgN��/��Vr��5��P�=ciXg�>=W��~5�p�;����1:�B���&�7_�Q��Ϟ�^��K��ݧ�����C�����:�����7wt�:Uw��WS�R�ɿ	�/PK   �|�X	� .W /   images/cca7adb9-3a17-4e0c-97e4-0d979b0e08a4.png���?���?��*t <�H��F)�ӱ�ϕ���3�)	!)BH���ͬrJbif�Y��m����>�>�?�w��vQ+]��n���z��47��}��]�=��?��|'&�Y
<�6�m�xD�{����G��d���v��X[�<bhb����C ���@����?�P	|��֕�G�����a��vpk�\Κ��o�Ğ����#�N�y�.$��}�lЄ�ԃ!��5�cm-O���577�5#�-B��N���T��?��������B���\i�H}?ҿ��T�J���s_	�����x����M�j��5��.' p�o����|�m����7��I�%�S��nW��369��o��fF`ټx�ۅ5���ɷ��:�c;�N�n�;��c�P@�ɨP������;�b�+�.6�h��6l����]�_�e��U����Zy[&�K"1 �޽-�d�U�hT��wB@`�:�d���ܝ�!p�*�[����	�[K��B���b�������+n�۪�<{�joS�[_�]<��%}p����d��kw�=�w-���G��O���?���}�Z���fsc3g��pD�?���+�gD�J$5���+��-��d�;$��IQ:��/V|)D�d
��'�(]|{]����1��1�������zn {�wQ�q�wo��pF�֏-`���i���1���R���Xl���Dn���}�s��o�\:p��]�����������k{�/���������3�JǤ_j���.��z���q��5���c�e`�}󦴰�>����1���B�Îs�Tlo߮N00�t�έ3g�Ω���-|=qD"C��~��X���]ݧ�ާ�VW��K-�++K�)���`�0Ԧ,զs�>ɰ���?������(��={D��J2��-'RWu~�� 
n/p��#�ܹs�2"e?H�}+�&dg],wҶ��>F@�w��ָ�:h�ꪪ=�ҩ�?<z��|�`��fz�>LO�^ԯ�
<����p)M{W��5闯�Z��ts���)I����ٹ|�Q����6�����}��mIK�)�f�6��\<Ǝ��T�[H;V��8�$����|ODͼ���������O��+ӽR�**�>>����]���6N)�*3{��t�w]	�t1��_�׮�SR2��}o+-/���t����ƥ�ѕ��p�M����<}k������5%x{F8���G������T�$��Ur��1����Xc\�U
��:c])OHh�����Ǧ���˫���ӽ��<�*�|
�Y���ˇ�߿[��z2Àw�h��4�tt�Xm㻰]��_<z$Sn��������C���^�X�F^��6vve�(#��h[�5�X_ۉ�@�'O5��^+[����ր@�����Y�)�/�܂�,ufM�w//.>���UH�VR�ot���8w�d3��[DN0��B)<H׹���V���w��Bz��87�����I�	�������R��+���U
���F��8�Q��K�~�4�>�8�d��a��;7��eeyy��{��'��<Z&��i�&&�������KOOO��m�$͏YQ�tIK��[���MQ�/X���$3�������4˼�t1�"jڏ�k�K����)v�������ޥ;�	�,��#���L;�;Vi�nW��n0�Y�u�>���o��bkk�qU-�Q�dfn��o�&������di]8��<\��xKS�tNT�'��ڄ֕���X���7�2E������t��������kz�1�Is�;�� 
�k����Yq+�c���^���c4��C����:����	������2R������p�=;�
�vqH�h� Ӵ������B��b]�E�Z�L��7�I��*/r��ijj�bJm�Fп��z���;��T���m:H�&_�1H�m���������i/���NP* (?(Լ�������з���_�|��ȣK���כcys��f²C��z�HN�����$���=�t�J���ʲ�8B}����O��kĦR:b�5��9�lj|4�y�����iW|z���%�sl��dp�OII�ɯ_�,H-F���_��ִ�,*�0�(���tTE ��B{m���X�������\��w-=��ׁ��te��o:��4/k��oz��%tL$t=�J�Tq����UTظ q�����[A��D�z��e�Lnd]�'�]C�c�g�׵�W�-����@(TP8Mq����Ҭ]��'^=.�o�ľ[_,o�?�)��!)img��<p���#`����]��b] //)-Mjj�8�<�v��uGGǈ�[%+�YT��1i��v$�[s�g�ddk���1�[�	6 ��6�>�V��0HE&�'�������Fp*�k�����cO�)@���[�7�,+ g#Xx����d�A�U�F�:%�����SCO/w�>��F���'�_ \��Ci�9�࠯[��̱13��z�*a�E�%>�v�D�^���&ئ��Fe�ꢒR��L��/-,�~�k�|��ӆ�����.~:Jk��\f��+�ΫZ!�U`������9:��:k���/����i���<yr��|���"y"B��y�`� ��Y&�4*��p4�d'0�N���[�tm6jȥ���5�^O������j����ޟ�����o=�>�ho����iO/e�����{� ��ܸQ �-I�9P��ӥ.� ��AF��YOC��?�0�SZ����a�'kb.G+S�_}c�D��q���p@e�[Ӝ>܀0���1�z82�]�e��2�����Mw�I����g�R�66��q�AQ�{��8M�{jj\.-)QZ�R��shh��@v�aaa�G�7bb�2s�#���R��K���� b��#ll� /A������Weӭ�OK�g���=���Z$�(3��� W'JA�f��e�����v�����-��]��%].�b���XO�V���;�$c�%_��M,1p�;����?d��|U��xѫ�e�@\Vv��N!�CI�^VbɊ��І�˲��j�dR��p; �YnS#r�>;�����su�z����kh\)��cfa�f?Y�����:���z�[޸�(r�r��<PP�S��_����HF�+����??ֺawv֗Ei� Z7B��Ƽ~д�+ؗJ�f�nle.�
k�~�.�k5?ǖLbs�7$�{xx����9���Խ�M^RFf���W�t�fݧrF�mb�&P��������Ib����![ B����S��+<�JY`	�#6$�nr���'Ws��*���Z�]��G�x9�����{msSR����4|ר����#���-���ȝQ!oNN�KJI�ۿR�R\^��5�N$��4��h}��ek����L���Lru��J�?� ��K<�(6�ɉ����(#�� ȓ��l�rs��wK�4o}sι�փY��!.*:��g����!��^+��-�-�/|������7nH����Ӂ[ۺb���#��O��Ѱ�@���p�� s��q�C')%m�!Iy� c'@ڤ/1���C�#�#��Noݗ���;7eF	���;���	J���7��j�C_i�壡��k��V�}l��y�J��Rxf���f�j-��ۙ���B�+;QF{b�� j�_�dΠLId2z+���j{�h�D�a�a@�J���ܑ>N�m�>U���c��d�\���\�aҼ���ɓ�\��,�p�!=�	�ٙ9kc/���b#c ��`M��\�����X�`nmܭ
DN��E����
��WI�i �!��X���)��)��!��%�o7�V�|e_(��ÆD����셉����Y��n�:�}W�u�h�'i����!�%hk�m�.iʹ�~���F���n�&��������{�޵]�n~aa��/E�Ǝ��|nm�VS���
��b@����|����t�G7�a��t<���Nk�:�������l��f��=��rs�}H�` ��ad���}J���4)��Ap�:����l�kr��מM� 6c�T$�K�8N����/�R�O%%��L��o��m��/=����XT����A
ǎAfkw���sw���2�1��h�h楃*�!3�*��3����`8d���Î_��!�#t�)���l@<��:��T_ yj|�3�QNt�V�^�˗ޏ8�VC+� z	X��ҀB.�����Fr�Ǐ[�z2�B �<���I����"}��n�ΟG`�`�-���Ɍ�FJߤ\�Ǻ�c�n^0<Լ-u��Rǆ?�;�V@��$$�#抓etJ��!�U16�*,"�����z� ���/�1��]���uf��H�H�S5�	|lq��^7�-��#�|=<�o�`
��Y����qk����%�J�ʞ�+Tr�3O�\'+���-8�޺8�����}s~d*3��@��F�gn�}�^̲Ď�ԝ��� �Su�!�E�zK6�� у�_�l�(c�<%�`s�v|s/�)p����f���+�?�+�t����4*R+m�����
圪z�F�^:U���?8�E��^�5lI0� �����?�������X���C�Z_��>c�lR��%x,`@�k\�wL<p`���P����[�By��7�T�\����1'��󷇝�ը����
�ʳGS�d�JtO����#�B)��ϯ�'�!aQK��k��}�>(	�#?� �8�E�M��j�)"n��YX���(L�k��o�)^0�K�*�QC[�cN�D�Uj8Oh�a��d�,�����&$� �!Lk��g��5)y����+b�#ܽ靽F�#�ؑJ�����0r;W+�&>䢪�VT�^٥8�C&��T�����M�Z��>���j)YU��ైcȍ��D��Ĳ������͖��2`� 7TT��=ڟ���c;>'���:� -l΃X�j���T���V�8v����&ND` "EZ���K�P�R�(ۀ(�:̝j bV<2I�}�]�!�K��l8���׸!�������Lf(�^f/-��k��9is��d��+�� P�#�ue�����;ow�? djG�餥ͦ\����K���=;w ƾ� �ʣ{̬�O��f$&ʪ>�8Q���Ub>(E�-E�M� ���-T�������O�����'<�:��W�ʊ2Rl�1M��\:d��!�x�&���	�Z��'�|�d� 7y�kz���q4!W�4��c���ų�����\�!��#:W�U:�w�b��_0�.HO�DfN!.h}i�m&G����r�s.�g����\8������$���n�B�������I)�>��m�����p��8Ѳ���+ �MɃ�:{����S]�cX	l���h���>�q}�?�����;_}#�F|J�v�/ߐ��5�Z�x-4e�~���{�B9�)���J���`��)�7��y���􁍏v8���1 �e����'�\�+3�U�(��1�CX^��r��x�$�$L����d�F��󿗖6��}���X�/u%�:�3bk��<��+e��j�b�`�����+Z;9��C"&��$c\��]cc��"���lho_�Lǒ�
n��ZE�T4����������/��MՈ������j�/�����$���
��m uh�L5g��ھ�>�li�u�JE���VDc�9��u%)%tT]�l��b��k�*_h��Q/@&ϴVʊąnN��7 �����t�wyD S���a�[��~�-C�M����n����J�o��#P�)���!��"BC`P��O^:U���`�M+�̃.���c���>��M���I��<ѵ��Hfz�Kۡ'���t�)d��jΉ����A��e��\��vcW��B\��~�-�Y;�N?`��]��)����G, ��/ �gXp�uNن�cV��MM��)�%"e5��Q��3�_{��+��We����+q��o?�ْ+�c��}ȏ�'~����V�����ѹ�f,veӡ���2� �%�O�Ц!8,/�%z���S�CC�ru#
��--��J���T 4��K��n��>܃��)���^�u��s���\cf��V�T�c�Ui�z�YE:-RE�V`���0"<�J�S�N��r.\�r�)
���MK@. �-VJ�nb��>��Q���Dpf� e�jw7�^����pxC�^Tyw��w5C[y���ٙ+��i�O�I.�5�;w_��
!cX�(/�ExhI�����|�f6"�P���n�H���+6���y�	Di�Tv���@! xP��+_�Ph5.l������d�#cA+�LA���L�Sqy�~� ~��X�w�"))I	=�w���'�������J�/ǔ����2�?���^�"MK�ۨm�4��"�:�Z]"qm�H�K�5j+c��wx؟��-�b��va�<�/ hJؔ' C�r���1��2��G�hH��j��OV}��}�rz���o��$5��u���\S�8�geg����#��Xt�W�K��	�k����իo5���/�"\{"g�AAw T��ܰz/��dLv�F��&��iGM<s��,N�(���W�Z�k��PN����x�M�DC7�]W�����R�;yƽň�lZ��źwBk�yî攅�|��.�_Ӵ�q`}$�p����3�R�m[^�fy�����Ο'�[)�N��](�X)u���  ��-p�.��{M�[�-��E�����lc8M���7V��o�]R#�an�{gQ+ϸ/^�D7�ǻ/�s~�o��1��G\m��֊�h�+�HuE���M3k��_�������S֕"�\[��Y��Nȡ�c.uu��L���E'X�G�������6A��ɢ�;�}���qrqA�ՙ�3~Rth�;�0|F�Zu�KFcnE�S{���]]@%�Tf2T�Kq.ݨ���ϽA�R�*�c����cz-����5�be`��?~t>Vߐ�2�J�|�^��]�[�������Af_�(Q2��(5���}Ծ�l��H�м�?C/b6��2z������:�8����3dxN��ډq���2 �xi��UJc�tr"Tϩ�2������2�)� �E�J��S����6����`
�G��������k�����3?OY�t�j�抦Bdw!��C��4��Բ������*мҙ�0�w�uѷǾ�ZTcW/Z+-�RG)�0< bA2��Z��4����V��r�HAS/��t�gg}{��jnł�9yBV֎�߈�*w�uз��� %�T���J�Y�B(Vs��ڝ����J*�F��V*�Y��3�C�(|CcwW6��~��+�_�z�k�VO�p�8
N`�Ƣ���{B�pf[xF��������^��N��B���N�K�0�a�X8����e���T�`������L�b?ʂP�!�R�<%X��<����.��Z�C�Ѫ�KƧ��Ԣ����MN�_�������V�ǝ���;���]���	9i̚��宯�/���<7�?;`l���^�5�ٳ؁[�;�wJ&�i�g��V��6�?���N]�����vs���G:\���ON`".�cq��z*���<"����ʂטs(��W����6S֟�1N4,@��c��;�>q�8�FK��oC"V-U]��+�_R�qU���5�,2V���������Bs,�r�j�)a��a9����4��#�+
5�w��`���X��TF�Ye)H�8qC'<���)�A�h�B�p��1�$[�W-E�;>�@,.p��]yQս3_��[-N�m�l��5�
 ���c�s)@��o�����\��j��(��thX�{P]]�ǰziq����.✎�'ľ9��Ǩ�w���=ո\�4������0��5~)���!(���P"��� ���NQ��㧻*хV^����P�>q���v����B�̵�8<4Jr��������8���Ve�����d�]���5'G��wG]������\nN��]q5N�~��r?B?��[�iN7����P���!�x�M�~X� �t)<�#E����x�uAK�y@��0%�2~�����Jp��Ђ�v��3 py�C���u�S,��P*��̀�z��f��¤6l�1�$ALJR�eZCwzH �(��}ys�2�*��Ћ��4�mr���9��qx��!�'�s�+Ih����^���,�,LUY�Ĩ�
���ApMEeu��(�nm�4�iv]�����گ>��z��)ۼ�m�C����V����mYBv�z:x0�
5��l�x���`�8����%7�D���'�����b�]:����1��|����ȬB��^�����t�B��<���A�j{�Ys<�\�bBZ�$}^\�P�~<�"W�cK�Q���e|�bȥjk�N�^���v��%q��΋C<FJ�iu�Z�f�G#Vi�Hi��o���g�����P!�?<Y̎
`2C9l@���u?[hΕ��B�w9�@H6�_�vI����
��ؚw��k2=fN�S�L^�iTG�.�b��+��nh'@�[/9Q�lg:D&���K���d�?~¦�
�� �b/��K㸾�����Ƅ���kx�Fr�樴��^���H�Z��ɀ�U�w��C�Y\�t��_��H�����$��^2��1]��� ��N�kv���O�#��E��}����K��kE_��^�*FQ8�ۖð�B��A���
X]�B�$P�qf�'�����{�A`�����?`�D�Tb&���������>[К�T���U~�7����J�m'��ۣ�������?*nE��i�-�k4��6Of�t�G,�Aw�����,>y��R���g��/שMH' 69�g�oǈ����=��a���@"�-�/�eM"�  �H>�ҁ|�81d�����YK_Q�xl���9^��]D�F|�����jxf���_���0m��@ j�[��u�a�P�޽ �!��䮘�\�9��l�0b�;P���)++�؜��������2򸯱1Z�r,���ub�̢�K�*;�����^3U]�f�f�s���RnR:w��l��_���kZ�~��E�$i���Zo��Gl��>���5���%X8���C��&�RB�WվQ�����H�L�dW3b�~���#6W��EU"?���D�]����F�p��a�VsQ�0��fJ�r��#6�����QY��4S7��u=������O#r\'��8t���ANE@�o@ ��X�nT9��g�V甔n���q�#�U��l�E(sڬ��{�hRqy��!��*o,~pO��3)wxR���q��ƾX�q�x@���ʚ��d#R��l�}�I��4h�vƫj��V$����o�8�e��fz6h{iC�6���|j��:�u�=t+�%E� �+��7� �1��N�%`��A�;��B�������5����k��s!GGv=}�ɇ��=w��?��,�ݶ���Y�����u���X����wK~d���0Q�TuGp2��W�@7�PG"���C���T������l���`uu0`�F�_Cޓ�'���%�YV��{<��j�وM�%ɝSV�g�C �?�O]*l��3����J]��zzj?O������RCq��әE��2�V��Q*��Y���C�\��d�@ |���ɜ��u���8����Z��t\hYW̗c:�99��%g@YI�So0�Myl�f��@�p&�pW��N��C��MaQa%ɤs�����hG̽30��� ��������&�y׹=��0�Ò`{�� ��Iޘ^��1�'V�[S�p�5�㽦���zr��Z��K��M'TM~��+��C`�8�+Hd1#�����]a���<?����/BE@��>©�صpjk��������6a�q�𙹵��:?��R�.�O~m�i���E�O�.4P�S!�O���#{-�`��%Vx#��Xz�~w=�J}�>�e�>���$�j.���l�4���?���k�9�����Hh/�!fg#>���z?��^W��ܦ�ks�H�H-}��@�1�9����`f����h�6=]"�h`h�PT�ٲ���n�̇�����M�Y�t��][N�~;���l�A����~9�i��9���D�a����M��>�]>Ɏ�TN�m"Ph�S��јT���_�;�ĉ����O��X�LAa�Mz_9�7F�cyT�)_���ѽkq#��΀w;t�	|Sa�p4������H�	ޖZ��+����I���Rr��	i�؞����� ��?�#�|�@�zf��'���K�+��Ȓ��i��a3='��q_J�Z=��V���S�#
����À�1(���\�ZBwhp]Ya��Ւ��h�h��^�umL�B���!��|�9UQ�hQ���@�Їk��a3c�bW��o���P�����ݡ��Ǥ�vK F�K�x+H�;�B㉤���ƃ%~�T�'�e��kuz,GE��j�	5|x�F��q�,�"�9��ʊ��L����1`|��_ �����{����J��߿;?�j�:*Z�ܽ(~����@�0��"�ok�.~��x�#��a&�x�imkA|�����U�g(U�i{���f���l�Ro���*+)q �o{��2�y�Ȃ8���q��{6�`�N~_}Z�Kb)�-��%��c�J��ݰ� ��ϔ�`	M(����>�H�2;���p�+\j�/4C�*������k��^Z�@~&����N���E��xR�#(����v����=a)��Z^ZZ���-p��.@N��5����]L�K�������}͆�}�򡑊�nCo�e�uW/Z	�߅e4��l6'1������FS�.,),i�H���c����|ѳ*'�������cm�oN��sM������ �l���"����խ�
]Ot��W���kt��)z�L-� +��0Rxn�!r�^�]���s�zS�`�� ~���;cf/y�_)����o�ɨ��
E�R�5�m�o*��ُ���H�4� J�V�����"�B����� 4_K���y{^�-`�0�����[Do
�މQ�[Ҭ�?΢2��8y���2�y��-	��9�s�b���ݫ{Ӓ�sW`�q��ah�y����X��U��,Ĭ������Dⶸ�mW$�ߞ&D`T��݊�ee& ��y���n�S�f�I���Б��� ��	J�=,?��t�S �G4�?������?ה��RU��ҍ��[������&�V�il����@�֩�tq5�g�T�'37���Oť�si���Ј������4�Г�&ֶ��\]��:�`��w< ,Y*�ژ�ѡ��1���k�z��GqK%�?��~t�Qq�Z�!��q�#,6%\���F�u��u�n��n>т�����}m8y�}����h��������f��G3%O�I����K���W�/���W���KI���ih_*%�� �tv�ϒo����̈զ/G��gQ�/K����:A��V�C%x�	��-F�f)×F�C�&��,v赵BQ�������E��qἵ�Y�p�߽���N����'��[^�Cn2G��n߃�d��8xN+E�d2&��v���M��йՠ=7���T9���_��,��ܛw�z����I��
rT�
^*-���P}��WD)�25�D�#�w��1� I��PC.|"��^�jvÏ�Ȳ<���Kݗ��+#	]��x���^������o��6�����K8�����)՟�O�A���5�w���H0�����0�=wRD����eW�ȒZ-)��0I��@��c�n��I� ����}�p��&)����K��I�ژ�-�q��a=���(^�k�~Cs���tB�d�>*�x_/�7�0�{�#���0;�p3�~0# �c�n]��O	�=Ҽ����T��}���ѕ�D٨������G�XÎz
y�n፫ڮ��\�0���*��'��o�w���O�/i)\�^։�]B2�C>ϴ�Wp�$�Ы��"���X]��9'`�ϔ>��˸���[Ƥ��'���6�Ea}�X�.�,*�y[�D�x�͐%zx�r��|B�;��ޘ�h���q{�����}sQ�Ү`p�M��(�%��{�~0l#�}K����Ls��vJ�|��|�IZ�QD"�!��U��8d�n$Lwx���5z!̹W�w�������=s�n�M����vђl䇏r�]��o ʻ�q��<-��n���HC`�^K�m�&)^x��F�2W�muɇؤ���ĹN9�L�)$#�������>C�>�(�,��B�)Q�g ��^Q���b�X�W���r���/�(��Ib� ��wjo2�wk�_À_����h޻wo� �+�!��@&P*l�*`���[`�?'�T\Xl���TX�/|5��1
5����&j`Ӿ�V(q�a�q��TSթ'�&}x��
k�eV�����r̫���1���Y����.HZ����ւ=�a��t�ZP�������l�,+<_J�<�D����U(oL#�\���=	�݁�ty���o�� qC������L��KE�6��6Lx�"cax����Ԁ�<�>
5�Y].�;���*�~Ի���u���(�yX��1�xE��N5����P��Z�v�Q��HN2�b�&�BQϔ ����!�Ji�~3EV�n�[h�����t	
8�[d��-�J�`#l ���G�}�|JT"K O�j�\�׷��I$�c9m��-��h�6��\ʫ��#��xш��)MI�
��+.�����^��D�y5Trs9 ���U���&f5���`Sr�y�꯳%E��}��9�}y	6a�M����*.[��DgGH~Yy9D ���K���d�!��Q?�mhhk70~󘊫u��ӕ=]��Y�2�##,���|�8���v+q����A�_��*�ثg�L>�c�{l�C3����h�U@ �J��0,�c�����E.q��"�y(/��}�YXCM�Up��8~ˎ��۹���Z�<�{�QFp���t� ����M|�i%f�%��6{혛�ۍvIY�l��*����7�N�!F��0}����K0.�������P���`���%�R��tw(�v@A�eE���0�S.��~g�}�<�;��8!_�R
k��T����x�`��jO���Iss/1��8�}���BCC�O��W}b�m]2�+%�ߕW۸j�`o
���Lu/��{�/�r�� �����-BO��S�0������4@aq��ȃ�P���n�/�.P�v�J�%G){]��t�9Ev��cI��kG�4,����^��v�i�<�����Z[]�k�����Ԧ`��7F^O''z	hD����!�#�������m!����������2ΰq�;��ǧ4�'{�8=&@��K.>V��Um&ר	s�[la�?Iᭂ-{�N�Y?���ڽB���C[�B����>�|cM�'ѣ@�����8���M����Rǀtx;�A�%�ow���~͆ڙ����^~�_L�V���0(�U@�%�'p�G���0�	u�-:_9�h~Za8��!-c�)"̊���M�������:_��ԡ����Ü%�n=R���uQr�*;[�K� 4ԘU ]�g B�I��0�� ь�~ 1��o[�5�^j�F+Z������[���-�v�zm_��S�|˿H�����|�Mvv��U����?ߋY����u4����M��%h��cbaD��ڑa�i5�R��p!���_��a����(f� �-��4x��)6Dk���V��Y��3�*��	��T��v=}^0�o8��ĕ�W�s�@�Ghݼ�����",��X�0�3uq�s������AH�S��e���\�Ĺ�CCf_(W1�:���@R�7�/��`x��V��0��zv;��o�kR�WsO��5WZ���><�J��>�z���r���n�O��y�[��r��L{�U���={b�����;�cWՉD�c�'l���T����~$�eG榥5����7��ܛ�ca��L�Q/���3�'�<�|%J��y[: �!m��]�k�ڟ5��p�JwE"Ӷ�~�U%���γ�IѴ�%������8ٕm��suY*E�5_g��1��@"ZARD���K� n)���瀼J�
3jT����So��b�x�����NBW��f��_:M�u�����b�zQ����I��ƶ�G��n�@�P�M�܎�Kл�; ��c�NO�:ȟg7~��H����p��#.c���s�5WrC\�cε��U�T-¡1uiJ_����];�̨5rtۋ2I�/�l/ci���c�S�;���g�.kl�\d	��D����M��J+�Ax���ț�Q���x��T�{#g�#��-��&��@g�����ڄ�F�{Q�7J�(��-ۀ�����v�~]����d	F�z��9<�p��+8��-��3�Py]�y-���keRT����1�6��/d���;��@�3��A�I����떨{��;.tt�z�\���^�}*Wg?}�xus��FS��o�G�DNM��|����9�_���M���P��ܤбgZЉ����#���������,��4�.�ތ6Z�W�e>2����{�O��<<�ћw,d �u���&��9+�lT�Ċ2�C�g���J��}��e԰���)�/���<L��c6%6�E_O~�b�'�#�ѕX5ڰ8v��� ����he�PS�(�Mͫ����b�ͅ804�SK�&�Uf*%O7),�>�]���o�R����d��-l c�8$  ��{�`"��"�23}�����&�8'��5��
�Z8���b�2��'��U���j>���@�;��ݔ+x���bf��D�Tך��0��y��Gٴ�� �	.E����q2=�)3r�����B������ڍ��Y�r6m�V+p�g�b
x��(�xy8í��)��C�l ����$�aN�Q���o��&$��%��F?q�w��剏�Ii���96��"������%��:B��p��e�h��C���Nv��F4C1�iNZ����l�]�*�،��w��_������ūXa�-q>�2K��Џ��>�U�/�X)ѿ]ɳ����;'g&  �r�r757����Vg�O�j����E�8�):x�ݓYJ5���h�)���C£I<��� ~��t�K�6;�>8>�]O�&tW�pB�+7��/x�Co*��Z�M����Rx3=74MJ!9g�QD�%C � !Ee��\j�Ү'����)8M���#�;���8��ImZڈ�f�@��ߌ��\�rBB��� �nȢ��怮=�İGU&��E�6���jg�ż�R -�I]I�fn�?Rc�-�1��Z�l���N	����f�[�$�x�^����z��������J�@̞}����q���4�:`FIX2+$��0�M�W�hs��ql�����Ʃ=u �ۨ�g:֗k�x|�:�8)%���3�tm�g�,  ������ϣǎ��h�6�y�v��z�"�]y�eł鋓��T�~BW��.�vU2|`^ף68k��������M�����Os5���)���	ăM�[������Y�P�7����*�4����(��b�\od�C9�Gt{i���j�|+`-���P^^�9��~������C�Z��N˳ ���y��N�QpMp�����ֆv�D�ė�y�q����P���ugD=j8�&L'�W��G	�m8^=Y�N-���`gE�J���Un���Q7";�jDv�P���	�:����1@���Q	wR�G��4�9��bq2��(�T�jBQϸ��j��z}N��d�/scܷˀ�Z����6Nt�j���IffJ)����.􋏅�,Y�%\�1.�s���H$�v!�2ЯIɇ�&a�]��,�@���i 0rX�=;`��mL��'H_�h�̘g��i�iV�k�ϨZS�e����\^A��vg-o�
pi��HJoJ��z���$��k۬����z"�}1�2���W�:�B�H�Mq�X�T��v�����e�����}.Z�ݹS�xM������u63py��.::Q%z�{P���Աj*K�J��m�U��@�zm�c	#ɔ��o󟢛�����{�we�mL�:]���8(�������#՝�9�H��
�k��C���2��;�B��7�6o����&����̉Z��f�d1��J���O �����
XZ�E���@���R�R���}y�4�#��xV:q�'J�b�:�(%lV�Y�Ɇ?�?6-�q�!#a!nB
�͌�\�֡_52��78@'*].�S pI���c� �*��s�0���U~a�t4[�y�t��I���%��lRz�.��r��X��L5�ڒO�����(4�^eeJ�q��@��!�~Q)u͟>~�t	��F9�p��'�־���Ͷ�&��`��ڼ!������2�� �pk�0N�4��2�>�7et��$%lmQ���3����߾�e�Z[qi���۵�=b=,���8���`S�{���Qܾl
��5���5��&�hHtlS8�{a^<��u�{�)�~��k�����[K���J�Rܓ�o�sf	7$�����Di�9w
٠��1M�.��0��u@�N�u�8��y��m�����ɴ�K��Ro������. {�K�xۺA{�^kϧ�c;H[����`E�?�������C֪C6H��Y-<��ʿ�ĩ�B�[;W��F�/>���o�`�c�a��j�_O4?Z�$����r���,����%�۾��[7�K
?p��D����G�K��?��h9G�t�����f�������a�B�N�ם6��[��E��z�o�"u�Ț�('���\2��**�z8~Ű�p}n����l݁P�o�Y�$���do*�"󄲝y�YY�J�����=���g�ᜳ��s�?���������<��y���󞀜F�ZA~����$�^V�Aޙ!/?~MN�B{��M��>�I7D����g�/�B���c��~J�-(�����%��b��j�p5Wܚ���N��+��(��U�%�_��Lf<�/��
|'1��:����"J�� ���xԵ���g㚺�}3���� ���m~ F���3q�AlL�>�룈q�s:*��"��5	���v��r��=@F�s��g���o��N�r^>41���'>����6�u��d���0���
�>�)1��u�~;�&��G�B;�.�Ԅ�~}�:���X�}@t�%����M�n��qH�(~`�����-ȧ��2iF�����D�Qٵ+LJk^�v��p��.V͇gB����������r�'r�R�����K�pQ����ߪ�f/�FW�%�#��b���=/�����v��p�=�*%J�d����]��2V�(WyR{~W���7ySH���zÓ$�oG�zk':,�.C�"-�<U;3�&m D��'��	�ʋsF�xm�����O�6��8�)`2%'��j1ؗ=Ra)pW%�{��񦔴��z_���H���fz���-)����0psêV����?~�x�|�ό�`Z�p�Y�u��:\�� 3k@2Z?����'"�䧇���L!e��H�/l
.�*��� ����N7d	��qf��T�������n"����Y�)|�l���h����N����{M�C'.c�$��FY��Ū�����	���Y�SR�i>C��x�Q��9�ʿ�Y81��x�C��8?;WN;��_��������8���}�dE�� Ι1`����ҫ4�'\���-����q�/8������?���B�D����\����C-�K�Ђ@P�oc�ĕ�t�#�:�IX���LA�~��n�;i���
ظ=�uս]Ǻl��
�,�M5X�Ab�<$��&�8�8&
 ����i�����djCg�F�tI����/Ǜ�Y��7fv�>U ֫�g���w�)��߯��`Ѵ����X�@��~_�=X{�`�տ2g���Rk�gZ�����%� ��5�δ�VX2u����`[ {�[H�<S��R�7��L�����%�.0����!�6<Y���ĳ���&Rd���Q��ޖ�_a�uЗVV��l��Ϣ�q�����[�'GY��ܰУ�$�M�H���[��:5��i�SXSG������[���{�`Q�m%�:�R@�.:��OrC<'b��� ,Ac��ØW"s��iIp�G3Sn��d"T�Szz��_�^n�/�,�\�`����A�u�~��)�K=�f���q�9��:0��
Dp�h@���]��¥�]�k�����ӓ�T2��K���F�hݸ����x�㇯����K�&��:is�'����b�#�cN���@B�ʞN����n����Xz�d�����hg󹍠�߄�T:��|B�{!� .>Q��f��*1�y_�"�p0c�~�ԗ! [�&}����9�/sT�I41�N��`8X߰�vq�����h��#d�n��ׯ��C���G|�M=�Bg�w^?_��'�S��Y�ӷg7�owg�6�R��1	}�U��>�=�c=F��t�K��ޙ�k@(��r��1�B�7�)�Sd���ZL�v�"I�|�Y��x���JV��g��ƫ���,����!�J�y�N$�N�څ.'Bk�Y�s�쟪8��tb��)n$.K$������=g!�g��R��ҧ+�T���:E�=E���������m�C%����
���ץ k�{��w���e�n�q�qݿ���;����.�����/���a$S%ɂ���s@��A��݊շ֥?svp:���� �c��'�&f�,��^_��vn-���9�R���밮���C�2ȴj�N�]c}�pP>��Ÿ�Q�w�Oۯx�hH8d�|E@�xY��R�o���8X��A�Uv����F�B�y��_���2`
*��K���g�hP*�d�E�h�e�(�U�We�w�=d;3[�UJ��[\@���.P�wP�V>E��*K�˯�b�n�d,����no��¾
�+��uR1N\�_� �2�{�I��Y��&���b��C�3Qhp�̡����	��3��|؉rvs��x���=�證3O�t8|~ͭ�[%�hG�-����@<���n���\@�������5���ye��!|l�����Q��\<��EZ��ƪ���[zKA3��]���ڪ�רgʊ����^4{�Y�H�h�-�w2SM��>3��ȝ�-���uqXҦ���xvxJKJ��&��X�����c (.-݀ �π�%��?K�u�$B]}�A��x�
��I�.�{��E��8 �nqPx����+�����+�	x�٧kCz�,�_�L�W&���l�H]����cm�6>�a�8<T)QE��/�`F#��1MZ���ls���[���W�޷AUP�v�qf�nЌ�.m˧���!x��"Ӳ_vV��x^^�|�?w���8E81�%�r:�wUkz]��<T1\c6 H_��@Pm�u�W_W���$U��*��;��#jآ�g�gb�����WXp(9���v���ב�3�{_t�ޛw?���{�����]²u�Kvk^�e�oY��y�f�f�|��U��������K(�L, WHQ�)�4���vK�A璡G���?y�^�yc�����A�-�uyl)h%|>���^�H9q\?��|�,�?���-�^�E�� ��.+w��GBk;���U��-ڜ�U=Y�>B#�<W�ظC���h�9$A����:���ς���|�J�����i����2d��[����H&��GU:�7�Jh���o�	X�}�0fܓI1e77�7�m�w��i�� ş�P�W�����w�Z�	34mRs�S��7��k.ٍ�;�%O*�q�HkP���*�cdD�Q�t��f�h���9��ܜm�,��/�B�>==�`��O�K�AI~v`.ds�����]��P��eFV��������{�c�������x���-Ȫ؁a�nW�nX��^w$�;�L6����.Z���}�%[����Q�)i0�{s3^�3�w���-�)n���`g�[����7�����D�&�$�W&���vE������A?��}�5,.�D0�ӫņ��*���Đ�"|�ˑ)l���W��	������}{B4���t�V���R���`���^���5z����A2��B�
It.��6��k�_�RvVW0�w���!Ju�����S�� p.:X_%v�\�3[Â���JD�XxAv즈��U�pw�L%-0IR�o��!���oo��S%%Ô;��K3]����F��l9��ڝ��~�	j�|�>�ڄ��'�����w��u>�FX�p���fַ�Oa�Liv�2!���r�<�៟j(_jZVܖ�Z������J�
~�t�/b6.��^�l��n>cB�(H��w�oO;d-v�Ịˠ]��D���s���8<dϓZQ�I��� 6�����Ȯ�*q���m T����Y)ހ
���1:&�~1�E��;����t��`;�_V�;)�)2L�P�x�9�%�v�+B�cm?PN�������1 �ݢɑ�|��5LM��fK eqD�ԓćyn�RR�a�
��U��ِ+�ܬa�޿$L�T$��#b��7� $e��c��Mx�	� �<���L/��}�B����O�G��+*��׺�BO�M��]�)P�u3y��[
D�4-�Z�g�V6T����������dL���zX��,���� S��<��Q3y<���'�'��e��I��#�ߏ;��JH�H�	�C� �9�����v��X�ټ��Ds^��q��q-z��o�-���Ar���c�u�����䄅{3[��?:Q��j(5m2w�ޞ���Y�����A�����?��4�e��ov"��g*	��U�1.��3�ޏ���l��(m��g#�i0��֕���aM��Ԩ��]AQ1v��5������&j�R��B�/��;<�Z�l�|WӾ	0�|y���	�c�L	MM����F'��ߧ����*��2X;sh=���*������"�Y[������Oi	v���e';�C�^��'G(�����ph���s����[�i��p�(��J�eӲ;g��AY��u�F6a`%�%�*3�-����m���K`�.5ȒށD� �~_.�S9I^�����L���Q��b���%��0.|�O�-_20���;1|�b����?:#b�H�T�f[=X:Q���3en|?"��B
���X��)puR����*���-2��t��g�8�IP���߼ڴ��ay�C�y|jw�QoG�n�}>���� 4��G5t�]�4�'�^F5�����%�I4��g�(T�)��n��@p�V1�%u3�����5b����=ɏ�~�y��w߭)�^�|���-wNE��7x�z�'╺��Qr�E������]o)���P]э�i6�G_%˸���֫��[僮��y��Uj�sfgU�k�!Ł��GQ��ͺJ��6i�x�'���0xz�M�7�!���	o��oww^�;���^�Ų�`f��qa�<P=�R�v��z.NI6tq��8��i.�߄F���2��c/���y�6��I#��ԗ�IkJ���˭�Յ�I��?iT�n$��[Pmh�AhR�\m�^�4�X�2SvR��:f��P�����W���V4ٰ�3=9"�r�D�(!C�������f:����!7+}��0er��=�)@W���%�7���/�6�Y��bL�5��e���V��<�C�B� �Z^�_U��Iɑv��ĥd��δ�v��C�J��$�rI�?� �������*R�lEe}$nΏ��dz8e��F�2Uϓ��re6)����G�h}�;/��(��$�0���B�K� vH@,���2=&C���r�z�:���/oo&o��ɱ��H����-�N�!F�?�g��j��un��Z�.��Ucd�Q�׷�1e͖<����(���.3��{�y�}����A�\6�(���B;�ۥ7u,%�/��c뭼u�b�����K�ͣ�ff],��8dhh��0�h�7�d�e�ޥ��e�yo�Yw�Z��q�B�0Г�hp���3�}����@Q{^SGk-��+h�$.X��[ U;�lk��Ԭ��T���$<I�ă�i��7S�R����Uˌ�Zr���7j�I��ST(y�D�wD�j�~P��jz��jr�V�M``��_�)�.�+WA���]��x������ix����|���ޗ ��=�H�}n�n�a��c���^������7��y��N�P�f�и�;�~φ5�#�U�q5cS���qM5d��&��}w��
҄4����3v��Kw�j~����|��$�&*��<�m��{B�ᆕ1}E��섔��V2v�����ZS�q��=)�X65B_E֚w׈%��p����K���B�V�2�����fi��$�H���4�'�m�N�Γ�v$���Q��POB�9�_��{m1���yJ
��_�P��$)�\�'���L�\��(&�ӝ�}����r�̀��#&�4��i�.�Q�!�Q�;����5A�y ؁� G��O<v`�������`�t�L�M1��TD9�I�7�oEف>����PݝK�|����	�L�iH�Aրy�v�lL	�ş6\��B����Z!ƨ.��fkJ�����U�}ZCW�(e�����x;ݏF�7I���<����k�����4�}�ib�����/;���|2� w�YU�~/� {\J�%�xN[�Q[�6S��[mL�21d~��:��Y:|
Y<�3�P2u�4�Q��B�&�#�ج�w���nX ;�>�X:�cUX��ua��"��q�R��q�9_z���˓K�{?�6�!*T<v[��K��M�q�%%���HP���m�'喢B��~��z��qu����Ө/_8����ؖ�p��,��؜�����������iO����څB�̮I78g8F���G��qZ��������?>�V�(m�$UK��C��P��^M�n�4����O?�k2�,��S��s��rgM�k�������G��~�&�y���N< �G��Rl���wSC]Jc�A���T8C��r^�9i7��I�-�y$!x�zg�<���^'jH�[�u�ϻ胼�_��y�{�k��@{�O�Xȿ��f��� ��4�r��`.0�soV�0q�5YĴi��b��5|�#;T�
�|�<��W#�����4#�y��ܰ�˨�j�*��MZ��K�v��'�Xm�i��.d��홟l���N����{?b'�@0�S>Y��3Z�X�bE��y!��?��Fh
R�Ѝ�7$����=�A��3��]���J|P}��MG�F}}���w��(���IRzK�ГԽW�~�p�?g�=8=r8ڇ����\�6��mNCX���{��A���������d�M�e
�{������B��R�[1@W�/��|p��Z�"���?j�Yd����%���f��̋QKm'$�h�JB@���n��tb�b�Z�+Bi���[���"%�3T�.��u���}�$���*&�7���h[���?��ϲ�7p��U�a�s�����ZnYc���0o�R�����:aB��]� T����X�U�WT�O�����;�m$��l����H�N�~������+6ځ��.G�ж����f����]ώ�f+H��l�� ���_߲�RZ�v��X�C��u����m�Rl��G���6t��	���=����6
�j�#���u�'���,�/|� LIW0��M%��j�b&1�g��6��)�2WY*��A���w��/T\׆�Q%�AlGY(�N~҂���ҽ�x=d�F���_�x�d*�g��M�9�-xA�O����'@"@��>l"�,�V���L��Va�Nۿj�����]m�������ȍ��Ɩ	Ɲ�Wr[��d�qM���^E�ܚ�z?��h�D�Ί@�nu���A4&ˢ�ꦄ�&!���e�K%%敗�F�dU(B-�ԥ�-����d��v	^���{�1m殼��
r��w�*�E����ü�TRRR���ӄ�4������>�a&�|�p����R��aIq�|Tj��Y���.�(/�lu�e��j��gW�%�O3(ޘ�� �P�7Ƞ�K@b�,���V�u!����,���un���U�Z�-�T60nȵ<5����G��M*���xw�)���~�5��k�����!��|��炨��{�����#���Iߏ!
�;n�+�ʎ���_\d��u�k���+����y9_n9E��-�L�����]�=_��q^x�/�9���$���#���]��MD� �4��fY�$V�*���5K��9�*�p<�LU��p��{�즹�'E-��H�dw1�{���6G>�x�-,�GN�"�	Y��P��*���$?�����ۄGH��$"Zʭ@Uc����Mí���9���|W�%��N�*{��{����1����r�ъ<��F�۟���7���Y��漻�T���c�cGGJI|�q����)ˁ�!�A��0L�Ou�:���!�M�/j���ͮ���K��*�n�$�w��~�]�Y�E{��ɵ��l�Kf�t�L�v4O&a�F���t�rlL%(��L�g�:�kJ�i˲�TnB1��U�H�!I�f�5�Ĳ��>-(8��9��D3��pf辙~@jꞢ����bZ��]���� K�Y����j�7�K���l\�^BXl�<�:?�܄N`������!��P��D�@������ڗ-�]��l��7�(;�C^5ӈ���jt�:ZƮ�P~I����;��I�]V	AZ7��-�:��A�%t�n[��Pꇩ��K�U�4����o)\���z՛�2$��px�d}�1���Qt�w��i�RvS�;�����ëqgj�2�Y-�ʘ����X_j�f1B�޲�̭ �0 BN��-��h���T�o;���~��~{���C��ǌ��7�x���%0���K_�����-3�N]_�tr�ٞۍ������P��%b����V�~�Ұ�R\J	�o���|JaT)�E�nSFc�.Áqp��.�H�Cr���H�NK��z�^��Ɠ�=����$Q�3E�+��n+�e�IC�f�
�����؁_Ơ�o�0?����p� ؀���Q1�O�/���0��������s�ų����>.���׉u�=��\!��_;8xoL5��G^BZ���9�����1��gW������t����>�>e����YM�A�JJ���1�W�@�҇_�����j�ꫝ��n�e�!�ٞR��V��\�
5�o�y���Ɖt������a�s�s&����
���	�?-ģ�hq�?k8�L�$�0_�Ů0G����Κ�.�F�BR���l������&�F⡿f�Wr�H��A��a��3�h	����
�z��ٴ��?�?�/��{wX9��t�T��I,�����5�n���ً}�Yf��+�/W��Z�6䦨ku�Z��ٍV�{�j"����a۪5��w2��YfJ��}[�c]�w��C��c�%�gh�~����G�;`����D�-I���IEZ;T`B��ؔ�ˁ��4x��6p�K7��E^`E���R ��~Q�\�#Yym鸟�g}�>�h4>;H 2���2��M�$f�u.�I�ܥ�Є��� ���1���/m�F%-n)՞��}������py�-~����VP�;mv�c�3��	�|v�l�٪��N%{ad��s���:��H���5���Wf�Bv 񋎗+���R'A�F����|덃0h��&��!�f�Ys������.�֚|
�Rw\�]���E���޺Q�ڨԡ�=t�?���n��I/Z�= �`�����B�L�c��A������6)������wk�6&�U�TN7����V7���f�u��+�:&�v��h���?���)��/�$?��T��e��_�7��-�(����\T��gC/ۏ%��k�����a�� �b�,�v#*{XX���9�	��I����v�D�A�5j��+�����n%?�T�V\��2zj����Ņ��;��*6R���
���+߽{�W&9n}�|�X���ms�s�m-��3DR�Ŵ`�:�,w��~�a�o��Zo����4�ޤ022�/�Vz]-��8�tj�j)���d�+����<f�N{��6��2ģ�5�RGO��<���KQ��C75Daۙn�
�s2�e��b�t���"ڛr�Q�a��yN~�e�N"����l?m ���q=����?Ϩ��|q�Q�j�����&dhڽ ���UK� �3��1���J���|x�����h��8�i������¤�K-���@����z��%G��Ŵ~��������Ų��)Pxl/=���5E���E<Z��(R�/��7y\:|�D�$�S�R	QԐ����%����<��P��ȼ5W���ˆ|@� ߊ�P��(µ.�dĜj�H���6!Z�g����,-�]���v�-�M�yC��$a�>�(�%}��J�/�" "$�/��K���%��3:ޙ�kz�r��݄�IH�6n����+�Ɯ��\D�"�Z*�"P3�ꠖD�#lŚW�� ��i7!k�P&����=B3�Ů;��Z�z&���U��Oi��������6���O�����3�1��e�Ջ���K�G�R|�iC�zY����DHӺ�����<���6�_�3�͜e�Ot��FTޑYr�?�᥼j5AW���6!+�P6��|��i8�q�����3G����˿gm�F��ڣW[�}�W,����~,B��`�;ލ��b�M��.uQ	��z�!I�J�U��>��b��b���d��L�-�X\�w�����F�q�Zٽ�*TQ��a��#h�8�=� ���dش��@Px;�E���c�hU�M�eB�����M#݌iDtvU�F��7���PZڔ4U�.Gn���A��HA�#7��Ko�����Y�d�|�wX�X�z�v=ݮ�(E�����X����)m���u��>��Ekv����+���ZMM������ˊ�2���lS<!<� �ˈ}�����ђ�4��40}1�C|��SW�Z������V��sAa�Jbh3I������S�pMcBz6g?qo9�U���M�_�s���i��!���W�@^c�5wk��x�덃]48� ȷ���)���ҡ^��xD�K�ܨM���p��!Ğ,����3x�[��ݟ7B�?7��[1�w&?��������G�WD���a.f����o���u%=��&�9�4y�^!����B~�\�|+/wg"J��!O>T7�j�k�,���5����1]p���Z*RQ_v>5��������͓��_��痣M�Uƫe�C���s������v�S�`�>6��J�)�$."�pc�+5W!��q�~&�S�����G��3��4˵���\h�c.t�q=٥\�8C�ͫI�E��'��}�%��	)2������Xz������˨~�1����[͵����
o[6�&\�-R��:Kx�K���ucͮ���v�!�%^0�F�ˇ�,�C��p�{�h�{��W� `}%o$���\X}�j�Q��q!�̮����*-��ݕ��|<�*�� ����F��k���������t7��2mZ�T����mNW��e&�� ��ӂ�Q<;eo0O敨�5jSnt�at��}eFx5��r�m�S����1�ݎ=�N?�c+�n��]��
&[t���������D�y�L�K����}�(O��VL]d��MY��*�VH��a�Lɒ��Vm�C
HH��GFbG�+��pje�n���Q��B�O�'t1V9x�O["�YB������?|Ƨ�(�Zd�P�TU�K�ջ�� _y�w��ܑ~�k8�iGN��fu�j����.L�Z�S�ah�*�nK�R��UM�_F���N�&k�	1B�����+E;��^!(���LJD�P��k!Ty�V_�q�].>���-�����l�W��#���`�J��?��]�r�1'��X`�ύe������ ��� �~�x�)t"���#�n׶��"J������-�|&��R_�OX��u.5�;��K�ֈ}���YOG�{�����f��G_��\)~â�t)���Ag���UO7k@�xX�,p�+�+�&�p9�j1�v曕������+S�h9~	u'Yc�����[����׶W^�Yot\�QL�ZKb������
b=�gk���;����п�p���b���*G%JB���	:F�VL1�S�o��/¥�
��څ�m��������6ۗ��]IC+����6�aZo�S�Z5AH�����fA��R�y�k/�6�[}��r�
�2^��˒�k�#w�	ǭHI&�g9c���4�	zv�g�{6ϳ<�q���'̷T�B��֗/%6fOq��ٸV �z&aX��]�𴫍��lꪔ�I�F��߼M�]A��y�&�U�jE70�"r>��)����u����x,���S[��g��X��OV1��G�7�k��+�.8mҊrQi" �V�(��J����S�����Ѥ������ڙ����E�"\zض�ޕ������������H��캪W�d����ֻ���&<s�fd�40��}�C�ᇌ�0�������3�RX��/K#�K���A�ۮ ��|͖b�[!.��|�ZU�H|��Wf�q$�U���<9pc\V�ۯ]m��>iߍ���e�;�m�-9�����V{9$,���ɓ^�B�Y*���]����W��n��{����v�CDpZs}gz�H-|���T`J����w���V@���(��N��,���jo��:�BE�L'�^]�����L���
�-�>4�iZ�"��_�-4ω2Ly=G-��{,[��c<�Űl7ĕ��� Z{		��v�4d��d��t�?����yף�!�OP١��(Lad��pv6\|�3;�\|�e|��1;*�-jX���&�0�\T5A�8�iEۊq8���ę�x�Ih�h���d��y�x��e�o�ˬ��9῎γ�;���J~�}�9��-�2h$f���.����7���	W��M�jZ�`-RV7��e��ٴے�l�5�O��AI6�K�)n�R`��h�V�@��9�����.�"6|4�0�ܗ�ON}ۼ�B.$�2j�<���4�\���h~�����eQ��R��ǟo��0r̔�Y��=��;%�v���y+���QK��
��5���A�{�����Y{>q	|j<&1��6�!p���lO���,5��[��p�N�ǫ�t~���7��wY�C��X��:�k��*�h���ߘ@jNl����ƀ�2⅃5���`����a���.m��=���'5�m���K� 	{5������I���.��z./~��I�Mt��\d{(����=�<��[+��������O��r�F,p�[CC%�q9����O��M�J�)�'X�Q���#4� 	���6��E,%��Xcq~?	�Ά�a�Dz�v'���v51��p�z1��������TD&QҲ�?��e�0�	J��q�	�Jv(:���K��]j�Ĥ�c�A�Q�0�l��u�{�v���f�V�_xJ�i"���������SOZe'�iܽ1�dJ��dH)��;�n����9)��d��'��,��!�_`K�a_�� �԰SA%�ي�C(zC.��:E����}f�嶏v���Kc�i��>z�;�$�2�%��}n��dD]��5ف6����~�^X�&"x-$�����ć�/�)��ko�b�����g���J�0 jŚ�adfO�Y�MN?����)�5K��Wt�(I� ��z��(!�:�@*��~��̒b�hY1�;�MV:�8N.CM*�Wy	��讟s �����ᘧ�9�P��d>��X����x�"+���ֽ�h��Y�P[xS����_��O����O�X:p�����&��O�����k�<cf�;����p���aH�'���{0r�4V�F��S3���P4N�ey�^������'�4��M�R+F����k�,����_�k<l��/�?E�0����'L>���JW�U͒�6��� �����U���������{�|)Brފ��4w˓�������$\����'5w���K$�mnK����� ��ᖵym��|�D^�vME^>�|�4Yb�wQ�/�״�R�_������1E�<7r��ttu�4?gfZ�N�V�ɿ���1������Gޞ�_��X�;xos���	��0�=�®�C%z�����#s�鋎��w>(&}H������'�t.��)����Zr�C*͏dJQ>v'��1h���[J�Lm�w�˒&iD�G8?�ԑ��]��{d%MCܻ2X�����zB;��������[Y�N���bW�`�̊���4[��e�)Y[Vş���x��ٻն��,h����JIEh�A����P��POT�
U�JHr���"�G9NUX(���3��|�?��gQ�A��A��wT}��O��ْ�e�A�SФ��/�� 2����a"�NW[%V��f�^I��(�|�^q����/�iEyAؤ`x:�rÅ~4���&�6ۛ����� Y2 ;`]��vrf�����d��b���O��8�e;�h�B���$��<ԯ K.>���|�!�����M>�a5�����A�i������J�f����7��H�a�(������!���ag9���n��	z{^�~ɰ"�gP^���;0p#^~�H}c��iJ����nXy܃��{Fy�i�4 v�u��?��/���N����O[U�ͨ�'1Vv��4�Y}u��?�Ѝ���M~T�h��D���5�6��zi�1=s)� ���p�q�}��I���h=H�K�4���١�X�� ��ύ�J����WX�~� '��@[UDx�����:nZn�$|�A�{�hH�:a���s�璏��w���,�*;����l���׺�.��&I�/g�pѲ�o.�P�,k8�Y�JP�錄�V�@]��Ų��VK��T8G`e�&����oIs�X�'S:H��CzT�6	�Yg�[iZ�}Ƀz��0��2J1�H��!�ݮ��|���{S��=�v^*�a�XjN<�=��d?����F0��v��$ئX(����:�	|�6�9Q.���0�0UpD2�7�Tn�6����� ��:rnh��8��#�o*��&&�����V�gљ��c�.��F�([�kp���p���-b�<z����5U#�������e֑R����p>nO:�n����?;#!Rʛ��H�/�g�՗�lώ�ΪH��(��=�:������o~���H��~�v�U<f�}(3=��k�3���Q
��b������Y�1R6�c�HS�x.}5���٤�߬}��$�:;m�g��6򵆫�u��Q5?a�F#���Ԉ:�T��#҉��d��(v��U�Ǝ�G��#@��5��C��ʺ� S�ma�V7�0��8��i7�Z������_��-�+x`�׎\� Jv�eb��v%aR.$��b�����`�5��
)�71]HS�y�6�1��2��c�mY��}�p���V��*M+���r�Ԥ�Ν�oL+ɜv0��]�ᮋM��ev��_�w�n~�zJ�����p�̊5���OJ����J[�]��
R�L�X��" ���1�B�ѿM���@�_K��H{��ޓ������M�V���ns�k�`��[l�n�wȹ��i]��(�d.w�ne�-�Z`>�?��)
�L٘4��/��:��#�L������� �L��J�{�nU�*�(�T����Y`��㤨�gP��-]%0�U��.��m���c���hǃ3촡6�%��Vyp��{�썙��1XVOf��z� �Q��}O�5�K�����hl��À���g�աJ�8x�z�
ݧ��{�e��??="!�TO.��k{�C〡(ś�7M�q�+xd�xV�j��ߊ	�ʬ!�.K�ɍX�~/��������¥QV.#�����Wb+r6ז8�5¡WZ�3ydc/Z���.�(X,��K5U{�<�ACTq����d���7�_��J�xiC8�����e؆�R]wD;D�#�MLLD��4��!�r�U֯��J?vZT����b���y6�Ĺ�l`�MW4^"��������$�%O}Ƃ���O�\���߹���4��7�Wd3N�P��z���!�t,/�!�NM0�OM�_�Мowm�q+���8�`�*π� ^����!��G^Q8��O�j�eR���P�0��^��qԏ�l�l��G5اSL�0}�*>���֪��`�-�Pn�����4�r���0�Vs�
ߪ�@(�Ө3�
�%���*�]L�ܤ#���K���+��"�xh���oUֆ>��$Gb�I��8�CQQ�y<�]f��x�1�L0Qt97�9���/P�TzY]��ױ�$q������/1'�r��Z5���--��kٻǐ���ZpA�Z�������f�}�ֹ��|�xe=2��0R>�n'���L�J�4�^]Z�"�*�\���O�30��JΠh��A��U�Ț�P!���솄��IƮ�#͑f�G\�����c����qD��փ����Z��fll��/ʐ>�}�G����6���ϼ�Q	�.$��7�_�h	e�5ܪ�~g���;
x�A�0�dĭ�p����ˮe�oQ��O�FT��z��!�I�d�HGԆ0׆��k5��»��ՒdmT�c����6�E2ɻ[�A:��䟸]���Ipj�x����p�M��~�F��X���-e��N���rj�n�P�'w93���c��U���x̲�eD$�醊~^��a_��^y`���\��A�^C�տ���~eX�N_a����и%Sa����o� ��.��� )�5JB�X��o&��˄��jy���|��^��{LzWz4 ��C-����/\[� ��Y/����?����qO���w;�%�VMF{�G�٧��+�T��� 4�� jG0�1��(!g!{z�I�Ou�3��-�Tzt=w[�,ݯ���ފ�!,R�+��G���[��vW���Qs�L�1,i�;c�K�#s �|��?@MkP�Rͼ�"]��'��מ{q�1|��u��7́�$F��+#��q��v��9s�K�I�����p�3�ǫ}pp��/\�K �)Η��������	LZf��L:}�v�G/��n�����|N!{KqTt�o��j��В�3�	+em}Cu��A���\�L�&���~��R��`��+3�r~E��GL���:�����]�_��/E�7�%���pY��a@�P{�b�'�ц�m6�a;��Y����֐S4�L�Z�3�m�Zw��ܑ�hHH'���Qb��m�ͺa`u�@���W#�32�|Jo��sX6�9�3��&����ox��.�^Q�k5e���hkӤ�TVV�Qo���������t��H�4�Q��� �)��HKK��0b�(-9�F7l4��2}~��u��s�������{�p�#��ߦ+�(U�����c�������7���;�#v���"�1�Z��*�a���{�F� �d�`̵��=#vǇ����H�J�j�B<Y�!exWRA+6.��£^�IM3 ���L-�R��|�KP�n0v��6"���J����#��X�]�8%v己���_���󗫟C!͙m�c�ޕ-�Dԧ��,T�s�	%�DF&�K�*�a����m���۷o���z2�׸O,v�J�x�\�+8���d���bI�9�%��ըA9Zh���o}�|�AE�*����5q[�(\��٧����K��K�Hf���S{-�W�F�~��+}BEƗ�<�'�`8s8I:#tY�m��W�dO蔌F&�j) �K��|��s�`���������E��dw6��'j��؀�����-�?S����g��ͣp��s�{�,P�	X6\�hE����$e�_\\��qrO`���Ү #� �+�L�� CpG���_����
ؽ:_�m��[4�>d�:.��Ӣ{�:P��7��{s�+�i���w������"�.��z*��ruf� ��g̞p�P���U)[fm��l3�_Rޭ&	q �]T<*.
�K꒸T�S�}�����`���&YQ����g�$0�hW��EmK��.Ս�Ɩ��`�X�����;�B�D;I˞���/��o�vݓ[�I[��@�|H������������nU��x��"[�vڱ��G��eq��4���T�Q��������x��Nc>��Z����Z]���}@qR�/,��2�O�VQ�3'>G�s������U����G<4�IϠ�F�V�Q���@9�O2�^�
����D,�ns~�u �=]����U�5��9̛M���v`��'�b4��N�["t�GI��\���F:��ZM��5�&�ӏ�Q�@q���2�!r��6�7�ڋA��魮mytu�s��~{�w"�̡�ǆ�;Z a�Ƕ�򧤦��_2`�gg���2Xn�`r�G��6��}eY]Ґ���Qy�ʈ⧈�~g)�T�w���A�-�a��Go�%�,V���!�`�9�;��j���o��_��d�'^���s{f��Vx>�[����ݘ��7/TǛ�{3?���tǘ<�^����*W��PD(�Qh�y��Nq�xɶ!:99�ϸ��Y�R�;��eP���FGcsv��A0VT���J˷vq�wDFl�+J��4�h��T�Ⱥy�4�mI��1�|����,�*Ҟ�)aS�>���n�;0k{�~y�r2X��c�F~O���]oS�-O�$Rla��J���S���[��U�a�>ϝ�.g��}y��T&C||g?�r��M1�^�?V����h�
�P�Ø7�\��� ������?R1�I�ӟm��OV�>��82 *%��w���Ƌ_��D�u$��ſK7,�J���"E{��S%^|�>.�k���:���܀��:"Ո��ޜ*��'��&�A����?�0�̓�]6�S;�ÌE���|�*{�#$��=��K+��U�5�m����LMM�K�V��z}�~E�i[�	�/�.�H���V��e�ȧ*��6F���?���^�T�,x�
�x��X��v�.�u4��hK&7�G�p(F��;<���U��XryR\\T����H
q7��'���������(�>
f����K�X�֙�F�&���{�����k��_��ۺ _jJ	yﰈJ��ZmubM���U��	Ứ�޷���!ׅ,��
T��_XM�7��B�-�Y�/�����&^߇�K�,]Li���pה8��xح�m�l�����7��L�K�^0T�����N��J���\S�å1������ݙHB�;�Y�C�R{��#��b��W��E�@ҭ͓#��*RB�撡M�7�9#h�Yz�}��`3Ë�͆^m����<���Ȇ�M��73Э���� ���?C3'_���%�,>T\�Fܚ����ը����s�](��Ls�ײ�HI���cT$'.��������]Gb��MrQ�Y���'�?\������d���]�g�c��P��	
XIgf��.WDk{ɒ��*��7)�9���ڱ�Ǎ{�&�b�̟}}d�U8�����F�S�{�r�(:�H���N��UNށ&�p���.�ĺ�.��珕D�B޽���b�G�$���G��_NEZ�[uj�:P�V}�*�OC4�V�/��X�~��{�׸��AV�3:#R���\�$w[�c�����Xh�Ȧ͚+K~���2"o�d�7�G�N�����
���P̑�����ҿ��,��~$P�f�<(��ź;+׎�1��1�5dd�-�%a�cL����ԛ�l�^�+l�N�Կ!-ґ��,
x2"���<DOk��P<=G�����]w��R�l�H���MP�Epտ^�w�o�D��~L^��-� ���(�
q8�ЩNF<p/c���7I=�w�g�TR��?M]zJ�@�ry����i.��ǏdLlҾ|yV>A�Q!�1�~�nfc4i'�.l�80C�+Lӵ�~5s'1��m�ΒHc9�R;���$9I��R�Qӥ�����|m�GkM-�����)0��Z{��}�����XCٜw�L�s�#��J�x�4�B��S���&8�����"�����]H��1��>�Y�=&s󲽳�s׃ʖ�c�P�5�w��ߍ���*���p��]��ȼ�6��F��Z<��e��@'[^�W-sX��IQ:�H�m�-�1�:\��hI6����ZS���yx\l4=�����AD����ň�J{�&9i��,C�T�N��Y���M�G��h;0�~�z����q�v��1m�,MV�h�0���n��. �J2}�i��J�~�Ƶ�mz�E���b��g�y������� �6�����D1P�@�?X��oگv��gs���c��j'�Xz�)��Lr��v��r���?r��	f�Hp�4��k1m�d��[��ݔ�%��g�q���>��w���,+-����66���J�5�m�~�f�#����w&�~�=�P���(K�YW�V��p��!���߁�����!�l�������,Y�zD?�p��Xg���.���5'��k��f��Go؁*�G�p��r��1�D��6���-v����˳����G�n�%�儖���	ut��,`ʼ;־6��=gX�@��!v�R*�,3^�7�?�_��S�w��
��6���F,���~Ӓ\5�c&5V� 2�<h�'�h����	�0��Z�p���heg�Hj']�G�u$����0W-!���km�1�V�C;�n��qN�?��K敀�?H��w;G{�/�\R�##L��yeIߖG#���,�X9�rP�NΕl�I��p���n�<G�He�E]��Vۯl���^��m��m��D�s7Mt�<�(���ݎBNG>R�y�\�R<�3ss5h^����>]:��9fu%�`J}��Y�j��ײ_�|�� <g
�`|���Ff2��H=�?���u}e��`R��E�6�{c����b�[6��^��2�=t\`H��v{U`�Gb����/[D�?��ٰ=���C���$�+r"g��|�s�Y�1b�c񎹄'Y���-G�TS�r��#�����5��>i[�����_�1Uw�Wγ���1V���.���O��Pk���:�wC��iB�o������nK�͍f�� �J'1qW�}�;Ki��		���6 D�V���,�EUi��B��W��Dg#?�gY�Q��b���|ǅ��I���R�w��� �ݎh�
‛��o6g����ԇ@1��r9�{���?�7��������4�K+h���ױ�k�܀ؔJֶ�{���Sa:����`��Z�����ԏ�}�I�f�;��M����C9��{������N(�T�yw�RoMc�n�^�߀L��`���꡽i�+��,�cvx��3�vD%��U�xs�y�o��OV���c����Q*l��_���M��K?������j�$����!���͞Gc���{y��y���Q~��9&!� �O�kV�Б䒏�M�`{)[�ȸ������˳`Y'J��9�q��B��;�GK��3}8�Ճ�Jf��ʕ@�ʊrpv:U��9x����Y�ٍ����l�~��
OQ��Տ@��@��u���{��-�Ey@�)\�$��~M%��'��'�2[ �����I�������r�ֽ��(�QR4p�c���۱�7j�������!�UUW�䰐V�)#U�{�b�� �������?VͰ��͋3>c߸��ܽ��$׷��;g3�zM��@���v�9�#���͚.}u�_Yc�9h|ܥB4F���~i�=� ��r�훓Hz��5��7�aC퓺���͜�U`�/'=��a�yQ�����/}`�v��f�uD���'�@�7+�U�
~�)8�GP�N[�X�����]��]滨e;\�/iQ
��������e�����څ3wŤ�.d���"�b�y��4Nkj/އ���m'�}���te�KZmm�-�v��{�7��T�T?�%YY�7�4��˦��zK�$޴�;V�Y�,;�_6���S�w֜�1w���"��]��ho�J_�����AIF��/�`�������}��\�Z%��|����3˿i<��q+y�dT^��7�_�ra���S�G����:�������x�v_���r�JMm����ˠ����[��n�gf��ۓ1���WS;����qq�9"��Y�:�M	V�I��s%�h'�<�Y�|%��1�3�
��0cWT\9g�B��EI�ʩ2��r�#�R����Ԫ�1"r�Q�JwG ӯ�X3�j�{�Ug�|c�7㍅ L�i.w~�Ȋ���.�K��P>n��߂Tt�'/�w��+-zc)0�zf������\��=I�:Aq�H���X��	%�� aE��F*�f����ٝ ����o|�7Pv�-���W�k�����o.�K�}�*�ҥ������J��饂,���A���8ertx��/�Z�������x*�QA����Qeg�b��A+[?�����9{��w����ǱG�3��4��⊿*k�q 'W�����ݪY$WH5��/^�@��$��<��Xɸ�,)bݬ���-m�||Yʎ]�#��Z)���3��x<��_y�ȑu4��ɐ/��<���\�G��Ÿ^j�.K�-�����É��p�"��r�6���~�ZZ���Y.,G��+�o��W����߁V�@o"����3\��)��&����Q[����@�Jܿom韲�R�V��*���`cK�hpV�Mܷ��aє	�D9hվ���]�5#h���[�g���cs�O��/�IkO ����X#.j�N�XLUAf⫏�Z��������U�/� �E.����1�/
ꅙeoJ�un��B���Z�lm���"�H1_�\��x����c�布��!+��a���9Q�љ@Ҧޔ
b�;\M���n��[NB/�ӻ	��?''�C��5qN��P��1�����%ʫ/�q+�}D�`������Y#H{O��N���6������HԸ�?޽Qʍ�L�(�'��o�ʦ!ګ<��G����k�3���$��Ժˡ�P�ֵgD��d�6�I��+f[֎J�H��0}�D���Dɟ�2�/K�tz'vR���������e�tk��ɘ{,�;a�}jXA$��z+Z �c���g���"�*��}.�@CakDfA93*��U�
�R��۵j��:��.U���c�U>�?
R�5tÞ\�%/�t�E��T���,�D��Ǻ����K=w
�|��\�Φ�:렋��m�˧Eu�❳�<����Ψ(�l�O"Y�M%�{������<�����S�}@�YH^�`��U��V��jZA�'j�/�����/��Lŀ�L-Je� >s*�fIZ�vQ[J	�zc�}��v�ƉwF}�$]=�h%�D�ז{2��#ZQH�Y���P"��	�,���_Ro�s.���G��S�ܮM����+�A=��3�8�9��ʸ�3c������yw\C2w��v�ڡ"��s�Q3�=~�h>鷷��?COೈ����>ssR@f���早(/�O�[�ҽ��4��l7��jT��5P{��	��կ=��6�l���Gt>�D�W=r9�*D�[kV%���{���,{5�OK!�*�[����&*�S��Zrׂ�2�1��Ax�t�x'����^�j��^�������󻦶6&�9�_NN^O��>.��Ǚb!�[=�%o�ZY������Y�j��=Y	�1�nT,��#��BL(�XvfM~I�8��ѕ������Q���dIu�m�Y��J�{�pYJN�>�c�׸s�r�ɭ]~���(��eUS��d	[��`��gdΦ�6��Ѧ�pi�9�T�P�i/sŵ�+m�W-C@��|��.�Ip	ZZ�\�Ѿ3�g������N�k�dgR�ΏH��(�vv�f"��G�[	���<�@�D,�����ji^�u��sW~�A=��L�w�+c�o1v9$���2q s�U��5�JT��p�&+��,�~����_^�9�߰zR9=�*��so>՝�XG�O`UbC\�凅���԰<�&�V�}r~�ȈB�n_����۵�w]L`���V�C����A�lYv�+�~>SX�������:�GP,�(7D�gvNY@b?j������5�~xؑ�8y�UcV��OP�3��ڼb��<��� �G�ċ��N��+�z�MH9j%�§D��&��o��Ɔ���rdWޟH��0�6o0t���ֱ�.1�U��x�~�qW�xbXC�ȭ�M��ӝ��0�KS��(��+���b��R&�Dv cC�:üKYI�J�4�Ɔ�G�^.�;7_�!_[%ά!]s��͘a����p�Ӄ����*�xX����LgͭR\#��q]d��4�EL�엛���8�9e�u���!�_m7g��y]��TX�iT���z#Jc�ڐ�J|��0��ab�=��鿸�id�G��g�{�Ɉ�����6�|45Xa�1��_����E�Z\T�~��c�����l��0#;˛�{�r�?��
��1|uԭ�����],�n;A�d��s)�(mz��Z��ݮ�H&����4;<[>M�Ǜ5�a1tWZʫX�0FI��;�7�a����X�澢K�����6��Y�<vRy��-����c8oxDi��d��r��	ԩ3���Q]�����_��pۖ��y󨰷\�^]D�Y�ړRK��k������<I�}�l���c��O����2n�YRǋ��!w�}�S�$W��])錹�~$������fds�eY�`3ʯ��P6^�`3=��Tv���-0��/��Ot��$�����C�2A�n̎�e�fc�2�O��[�z��ü�&�}��������e�l"jZ�����|�7�W���vϜ�ݶ����O��y@��Z֤�j�a�ҭ�4���}�BӞ!.�^́�c$�-u1rm�L��a�-��M2Tl����D����Ά�PK�Y|��`��}��s}�4Q�)�n���X��4JR�{��,ˁkX�F�MV���OB����1�]fcq�̰݇)���8s�ą�B4�u*��	�9�Ѳ
v3��ND)~a��B�m��̔�b��J�,��ϕ�rxHa��/j-_�����f�=d�-�O�QPz�E1��v�;�S[լٵn�iVl.���\騔!7P]�5�M&D��@.����i���|Ա}���z?�[����>�h�Wy`�a�W o��F�퍒۹������G"���{ȹ4g&��m�x�3�`��,1Rv�xb\�{^�
�q�|���6��F? ؈x�q���^���B>�=�b�l�`���v`�
�h��kaI�g��^��ܬ[b�)���!Ƿ����V�y�O���4�e���t`z_���,v6��0����E�S��Lߟ*�����D^��0��~��v�����x�:�Ju�|�VꅄЈCs����q�Sύ�%X�c�O+�汛ě�JH�1}��b=�����֌e%������{��q�״���]x�s/N썳��m���k��`�l}�ŝ,fM�\�>�vQ��u��8���7;�u��/?t��]K� ԝل��=C_�i�)���bC��_2qY$�5(��Xi��u_ ����J��d���k�8����PE92#C�G[���zV�C��ؤ�	�*�|�Ҡ�!�/�;�f�NÓ����֗��]���Mؙ��^e��2�����Z����x���!�|�`���Y����9�4{�SkH�l��۵6��*;5\A��(U5[i�k#�pL�_�/��kS����'�y��t�pOw��һ�

I��A�<w�����QU60u�!��^�z����f��d.Q�4�C��/9�flwj���(�I�ԾvXJ��2� @b=-���z�Dy���럭#��P���Y�M��ѕ֗?��>1}o�S�T��M[��"A����o�*|-0��i��&�,���Ա�Z]����;0ǂ<���^��QN]K3;uK����9�-�W�b��ʶ��StS��^����3�Y7^(���z�6 )4�TB����|l�J�K�z�5�M�_�{;���]��b�uL/g�}��6^�����gb�����ōk��u�Ɗ&�ū��pM��	5��ߛ^Yì�`;��[;��"���>���o�
;�:�,�����'�b��Iӥ{���i��Q���Y��0��h�p�l��u��Cy 	��+-e�} 	����mr�=>���|������,>���}9t�w�s$�����gN�zC��B�	R9�C�.d�|�c����������_�z#=�tΪ9�{��f@�To{�T��]�Ũ��H�n�ʕ�X�w�fOД��Vj���@�����BP>o>h!N�*�MC��_�j]З!��n� 7�Jx���F��~�j?+��	�g�X�۷�Ba;W�^ìo���5������%�k�y�(gBxKx�v9������Es������e�խ����'���_��ЈՑ�����YnLZ�!a��)�p�g�/���e��.\Iޗ�������G����Hf��S�J)���	 S�VT�O˂�zD�A��%�w�R��DQ�k��g����韞���;���]3�:Z�a�G��}�Έ|���͋��-d��J 3f6�1}�]we��_��m��C;to�.�@�U8泅�xSL�(źF�*��R�*��Ae=Ř?��\Sϧ����2%!L���e��8�����M���(A�k���1憬�eXhl2;��?y/y�m_���T���V��?�:|�58�
C�U�e��bgxe���}�8����NlPX�J��T��b#�m���-q>�0��#�ߑ��m�7�U���*���ao��o����!"sxkUJ�D��q���&�/�P�da���=�e���I�~�l�� ����J7]ȟ�C���Gۈ5pX�[�y}^��l�B/X?"�	��U��X�����UTW�d^�f���K�O[�7ʶ���u@A�vr��j�j4 7nJ����qUy�vn]�p����T�ˏP^�o�':O?G���TgͼyK�L�8%!��r��vV��'����o$�	��d�Z��h�S���I�G�0�~��PV���ٻT]z>4�j�������s��h�>%a��8�n)�lIt�(��7 ;�]��D�5�H�_q79�٭!\A˽���Gq:�l-vHQ�)�庲W~���%{��9��#���F��� (�ޛZUy�r(�@���(L2����)=��3^6"9��bi'���^���w��H34R-z��WY��2⺁�Y��]^eN4�Y������:�ds�-��W��q'�9�CuK(�o�����@���T�/�d�v����"=���ض!-z|�1~]���c(ݪ=��Jj"uF]p�T�Q�@�@��O��.P�gU~�%�N�Z?�ٗ=g����mF��,��]�Q������Ҵ�T�m��k��X>�ل�Ug�"R����i���#�o��|�<������Q['�;x�~ `�7����S���ƧT�s�aT�Nێ��=cU�;*�J�R��5��Bfq��@�X���%�K�� /�4wև�&Ԫ�WŴW�W��Y¤R����5������R�{�ٗ��N�|�e��r�Ά�߬��=�� E�?~C+�� �Z�Qh��$ek9��KBwx3YRwN�	&utm�!W�_�[��s�V�<e���S�}��5l�_)S,��ԩx ��
��Ok6����]�]~�D�|.�U��A]4z�����u����[�h|W����^�,�ԡ;��#0bD�#�i_5C��2�����]���6z�ypQ7���{̆�po�%�9�j��&�n�N�X?�'��e����x���Y��z_��`���z�WV!���yp����z��ox���%��۸Ise����s��(��tF�U�%3�ی��[���D\͘��B���A��00�Ռ��G^Ț��L�����O�d�fW�Y�ٲt����9'ã��I�`�[���r�����$��>G����T-����̩���P��)���נ
H��:�/��76���:W���8��U�n3s���HC����[�Ag���7�z���4xKԈ&���Uqz��� 䢏��U�>Tw�Қ��}D��&7�������z�����ג�s0��H>���&d��Iz�Ay�r۷�p|7���o:�2t��B�!��i��!�d���ϱ�T�ɗ�;�M����n�v�!O���9]�;��w|�����[}�CzF�S�x�b�m�?�� �t?id�3�pF�mz^�3����R�L%�:%@
c��H�9�O�O���Movff�5TL�:��p
�+�Jo��?��^Z����L�m;wn؉E�jI��<�!C}PI}��^)�෈���Ug+��LrK)|�֨��am����;���מ�='d% 4��*�ѼQZ:��b�SHY~+i3̋���+S��)Qm�����	Yc!�C��.�UV��C�t���B�d%'���DU�JS�m��k�V�_��>G�.[�z(V���m��	w��g��Hc����Ⱦ9���پ���֭���P�
�q+}^N�����9Oi�����w[�?����qFꮞ���j�aM��%vgT��]܂ǏzGx�'/[�:`��DO�(e�������v��d�"�~g�m,#A�K7lx�-�����S��S:Jۿ�nӓ�Ϩp����ޥ�ݳ�F����鼐���P�pݣ����[�����{��W�c�GR�l�E��a�=�iUlU<���o���B���mE��ىn�*�@2;`u�/<��9�����y�E�u�V���Y^���E��A�2$���?�?�<���J��z���'�^�B/�����i�xK//��J��h����H���"1��~�*+s�=�^��ʖ/G}M��M���wa�3u��J.���^���2^�2��IBv`yx|_��Om��D���3��>#�j:�7�I��_"ܛ���*�ɸ�v :���`�L]C#N/f�[_��L������fPD(��'����T�5��4Q��F8�
Ȅ���'��`K��+���W�g�P��[<�e�=.F�g-�v.�/�F^�=.̄�lz�p�+Y^R��*�x��]�����cAtC���`t�j����FP���^Q5\D�h�c��&q���b�^n}כ��;GQ��3Y�
�"��F��qN�BQ;�Hp�
b��7�9�����E�)��p�eFD�~��3�a0֓�[Q��L1���/���_�4�G(Ǯ$�ds#X؀#�	�d����N�b�����lL�V};��X��Ӝͪ5a�:�qx�������2O� �ɸ#��Rقq���I�OSI�u/�֨�J�`e���Z������`M��/M?#t�#�����;�Ch��c�
��;3���e���L�2���ć�7�|��o�_�*t��:�����{e$T29P�)!u����ݤ!aΑ}���욢Ѫ�%`<�����}��E���RN<ϹC���_J\I�-T��f�����Y�w&�R&�� �r:���?��'Y���ނ_�6Q��-Bn���.%Ltaٖ���0�G��R%�%V�31P�C��'�<�U9�T3X"����s��J�����Y�h>��I��Y"CI&���0|y�����41�맸һ]�YV�ʍ��Lg�V?�j� �֖8^�X"��F�:.fĶ�7�|��n-xy�_�O\�4Ol��y����E���ml�@5;�ڨ��K��	C5e`vЅo���M��^'߱�e��WÇu�ڭ��m�+?S�Mw�żՌ4JHH02�c�[I7�e?�S�35޻y�I�s8T�~%����Z9]���{�+��d@W��@�z��(��{��f�ĘN��\ �u�T����}@�]��ߺ(�u�W ���t-�����L|i{'eG������.t���4�R���Jm�e�I��Wh��M��L�ѿٍ�� !��Q��@.ͱK�V�Ҫ(P�60 �����~�2G z����O��x{����=g�C���'ŵ��fG]�BUv>g��B�=I�_wT2B�?�ѐNJ��6��	�1��������	)^�����}�P_^�j#I@ćmֵ �vI
Ⱦrvjʛ.R~���H�i�D�3�*�3����Q��ѹYa��G�������	��~x�Ñ^����"&�,���ČFRv�	����X���c�7!�:�9�m�	u��(�s��p1�����FJ3����w��uH���ܖyl���g���ו�[+B#(7�A�{�K�Yo�f5HB�H�����Q�q�#���U��-FY�k܊�}[���e��hgcY�8��b��Tt.�4��v��\mw����Ӎ��Yd}��k,�:7=UC "�-b${F�g�����7�.Ր�4�&1JUI��>%�=\�_{sX�E_G���[ivn΂���@���Ȩ����G�4��1&�{�3��H�m�
"�c=��]/DN�^1a9��7��Ѥs�	�"�JD�=��ow��^��V� �k��3*Ta�_�9ys�d�h����_���ВW��	���_8NIM���Ap���F��1B��&\D�����}�\���D����WѢ�GGݱ��J�n���	�w{�DA����S�� 揋P^�]�vu96ne��-.��et{�8gl����lMa6Gi=���D����7�'�2H�M(��N�_��h�O�1Ѕa	��)�Y!���mбdR�q��՛{�3e��jdA$Qs��b�d��>���*<�����ۮgV!U�oI�+r���'�A�
�'�x+��l��'�[n�Y[�+��z^�5��o*Wl�PJ]�m�����x�G`�O�%���k���n��Q;f��%v�����7��:,%�I�d�VhkR�qN\F��[�_y�z�0k�p���\�]�*�.���~�yƾQ ��ֶ��������X��
�����V5Jb��l7>S	�����=�SZa����@����ي���9��n�e+$�}�F�3�*B�_��<&s�͘�V*��v�����y��Z��u��e�(u�&~E�m�QR����/�$��~�$�L_R��	Dg4�k�Ng�`Eg��&�� M���91O)�6�;��6{W7��ߙI}�q������P��kc�ф;Gv'��̔����)>?�Ur�{>zf76b&x�xA4��Nk]��#6�u���~���a�m�){u˥�T����H�����f����'?{p�wC�B��c��� XI>�~v�Y�1 L>����0��|�חV3�S��B�"�,o�����(&�H��壖�it>��j<x�)�~~�Cr2���c|s�� o��H�C�K����Ry��\�2��J�
'i<�s6=����(�8�B5m��kd�T8S�c����y��u�)�$�Rʈ��L��M�r�w��{�S`5�+�j�؞��8�_z9�ѣ;���Y��`~��C��
M�כ����=��I��3^:j�#��܏4���g�@�*y�7�syOMx�e����3���t�9Ň��e(\�?��8B):oH�u�Ӄ^)b�׾>v�BJn�}�$ʅ0�U�0VIxWl�.FrJ��H���lS!+.�H/��L��c��r��o^6|�-/ȯ������*c��^,�\ZS���E$�犞CU�t�W��͆���>���暍���������4�z�MU���_/[��r�6)�n{�o�n��3z`:�#p$3.(p�%9�Z[w�V&dY�QhS~�a0�o�
@�t��Cz?��/~��o��Ah����l�S�sA�Ò����>)��^�-�<��ֈa�s��x��Qf�&�@�"<'u�%���n����#g�@|�S�&���_�3tO��Z>��Ӄ4]ZՋ�j�%��a����ߊ�8��鋀�MM?"���g��ŉ�h�W)No��Y((�X��������j��7�� �Y�s_{4�f�!N�^�/�Kq��[{\H1ڃk!�X�+aB!��N��:�l�<{��̑iPA[�0����@lX��ו~v��rE�/	��i~����1B����_k�lރu��gDx������6!�A��}�r��,.�~2:�f�E��U��5��H�T�a[���bW̅���C��t��R2��	g���J�G� ���xf$4h��픗�9�3���"LEkBl��Zf<������Ͼř<w��=� �#Ц�;�]�]�`Y���{i6���L���;�n��u�a�����	�a�S4�`�
�f�i��O���E�B�� -�a���s�cdc�<p�7vO$�{H�{.߳���v��J�t�p��S�^��ٜ%�l��ÔJ&�V�Ƹ<�C�h}���V	�N_�U�u���t`7����ˮ"���V��s}�R�����Q���ro�{�$K�m��{���4�ϩA���N�-��0tṸ�o^��Q��O+���6F�����`��z(���7�,����?ߣʃ��Z�ccI99;�� �骏�\]m��6-A�a� VG���W��Q�� ��/�o�᷼�ІTP�JW����J�(s�zJ9���P|�����"�ȓ����	�L��[K�2�oM��%��xS~�[�S�b�Qj&yy��K\xOn�i�{q��V��Y�	��G���>�B���+�GZi����ZwJ��{^R��d�͇���4�F��o��]��zV��dgߌ�����,;%�/l�i.�9��G,�s(K���ͽ*�a��p���a�r&)�����P���}�ptź���7�k��3�ؐ�M����o��he�,�\�給�y #k�x�JnZ���`�&��P�c�'le�����Xz�)4�f�ݼ���6����}��Զ�c'�aDѪ7"�(�	O���dEqڤ�xt�{���Z�}�0X;�K�Ng��GD�)B&0�)���I&�}:���J�ǳg��߁_�������+��'N��7�+)3b��^�GXSow�����z�:5/��?r�|G�?|}��-���~Uo~%�<��SdIUC�{P����AsO�ܵ�P���tr���<<'c�u��7����?���ﴹ��a�)�9�s����^?�r�L��>l�oߟG�:wRi��[w*�C��[�
���l�9��Qʟ���͟	��
@4���Q���z�^G�_C�wkS��Y�.�L�sK�ɿ�i�}���(�@�vupC�䆄8��ѷ�P8���~�^x���H�����	{�T��{��B]��!����u���!�Vh1��� �������'u��`(9������)���>���g]��%V���G��i(��� ��b�f~���$�����K_���ב��*���@�H(g���E����T6ml��BM -P·�9�(^��j�^���hN�2ҧ�����>Ǔ�D!#a�UYy�"�J�b���@KJy�Y�h!��k8Y1�y���J&�)��M�[h4
�{U��5���:j����D�����������" v�9ǯ|���oEz�HMOFK}玳���K3�us�nq'Cq6��1HH��N�	�=܎pY�mI���<�?}�]g���8��Yr�iؠ}��7d�������e���H	a�o�*]�J�	ˆ���8^���I������G>,Y�~����ﳹ&Gb��0�!T��@�@#-9:��~�Vw������/?���� #/[e�˄O�W<���R8[���nb����ǀp`�D�'W"�r�kq��>�lR�l��ѽz3?M�Z��ǖ��Yv����%��{ʦG��xm���Z|3Iw벋��6�;�;��n%�շ��6��ҥM��٪�M���h䆅`G�W
W��?��;�7��ޫj������tش�7���j�V	J��Z{��W��"f�;b�������/�9�s����{��}-BqWq�@t��s�#ё��Tl�>w'[�k�uW��$i��a��~��/�T�H�:���i�E/��?xĲ��9P��<q_ۮ9X9k ���ڢ����n8����[h_`���u��x���4�r�%Cw�rh�+�k�0��,��U �&�m��S���J��x�I�h���z��!����%R�Bw.p��}����s�)�Q oAy�� ���4�����*Fpi�a��d�}�Q�A�&��~��K��fԀ��u�ύJ�uؚV=X����ո^̼��F����%�H� ������j�C_���_x���PzF��7i�V���
U�1*��m4�hx�]2��<ь��I(�t1x��#[���2id�� ��]�o��ɮ��������A�n��#�Y���<��!(;b�oT��EU�|�y���H`����'vo��qNK��MȪ�Uu@��}j�u.A�,E[ߟ��s�oI���W�~��Ә�QZ���x�7��+M<>��@�Y��uZs����f֔jhy�����g2��ݾ���__��j'�G){0I������c`���#&��$J26���,=�Q7]�p�s��v b���>d�CA^�>���1^�r��ڞKs!�Z?M�������b�?v��5�9�7�5�
D��V|@l�ĈV�,��s0\��1x;}�~B!e#d�U���;���-Rnu��� ��,
�ˉ"5��Wn!q�.��`[�`���\x�����M��V���W|�����ٌ�(f�J#R��mE��,�H�l,�-j�\�R��C[��b��m��h?����7��.s�	�~p�o����Y��H�]+�	�<�c(�C�sW����pys��6@���U�Mn;��IM8f�e"W��|(�x�~t${�_�Ҏ2��*����.P�('��FT0zilo��d���\uC���
��;��Υ��4�4F��k��s�z����}~~ʅ�.CWϾӨ Rz7j7�(�j�!4`�両��VCG9͙�|�����3:7h����	Y\��t^����ja�7�H��?��^��9~��(�C���n���7R^�KFT�'ɦ�ʢV-�t�V����6��?Qc q>�ڜ�_�\J&,!��[^���X�u���b��A��a���(.s��GJ�M�k���Bf�G��z[��d*�F�`�����?] a��21r��Z��v�ƣ�A�9�JB�/ȑYk�4�]_B���?o?�m�|�*Qu�c��hM��#���4.��Nx�M�=�1j��G�d�iC>Nň}��w� ����ϻ3�ˆU�����>J��؝9}�����X9Ҽ���k�����r�~�����w@�+7�'������~�j0}�6��Ѣ姀1��������A�K��V�o�]`�n�.]���>sR#̨�48�^����3=~ŇZ�l�ȉFC��������-f�7���1��uE�+!f��=� �]��Ta ����~K�Z����r���?��X��W W�u'x��r%�&i�4k+Y'i{�Zo�(��Gm濪���ϭp���s�����@>��8=�P��w�]/.�������A��d���N�d\%�.!���d�8�;�cq��J],2��	�9t���
���.��[<
)~+{Y���#��-��J%}��g�������ʦޒU�C݈��V�x/	�,�t��n$��VΖb�C"^��T5W��5��Ԕ\u��aunr�umAǣ6X��b"V�����5.]�7���|ޱ������۟`��9AU�������G�D7$r���d)�\���I_��N��»�Q��p��d�@�	�lI��b��k/����w!��Ŏ:cά?�w�;an��ʐ�&@fc��@*��("M=dNz"�V�h.�������Q�ԕ"��C���dE&l�Ȫmӆ+�Np~�5�x'��X��'�_0��X-��ܯ��0���.ӻ��n�g�A������	����r�\��D��~��^����O,Y���3���Ӫs;I�0�Rk����h�t�0YTh��I�%I���h��5� A���U*���?�7t����@�j8��c	���U�w��E��t�
��S�Y)@|�3���	s>ɞD�`��c��>~��zY���=ោ��^ܸ��P��\k�� �������dW�������w½00�兢���.tܝf3欓�b_v*dhS��u��理O�Ф��3�1�g��~�iRE?���;��{j2�M49"�7֎cP�0���ϖ�"bde��.��B����?o��gA�i�)�h�z�/㾦*�o�µh��P�k��dJ���Dm�N���t�4&�N����'�}nr���Oq���UO���oc�����:���!�3|t`8���ډ�ꂏ��D׵Z0qS�,�<[���͓y��I��+�a�����I���h���r��8'��f�� 	�����ū�Q�X?`W�,�&6���Q=�Y���/֤� M6v��:@�8�qRv��Yq���m�<cۢ�Įr�b��)Lq�Y�Ԥ�����qx��hjյ�6R����}@7.�1^4���z��z��A��-�E.��1���m�8��%*���oރ����9P@����ω�{��;0�Y�;�c8��&\�U 	�d k���z��G���|�n�>��8.{�O��S���S6��'\w�e���"��37������~~��]�հ�B�2�0�Z��?ū��sx ��<�-����K�/�=U]WY���i+MV�-����h%9[Y�ż���i�$��#<5�I�6����&|�4����(�J�m�o`�'_�2]^0��1q�;�����B�U��\�3��>��$����H��x�]�&����x6F1����8Ϳ�&�9S�е����rz�2v?�
 �l�����2L�[GH��?�3�Ӄ+�qȷ5K�(�{�~,'2YݯPP7���)�xf~�M������0�\��)�����,!��68ԍ5���r)Y�����Üc5�5�J
ޜ�*M��z��{ߗ���ᾔ�F�c:o�J}@œ$`��vwux+�!M�����=��<���Ss�"�����f��%��TX��R� C�o�8���p�mNO�[*tbn����Bc8zt;>⏨�s�\�+dk}A�Ls��=m�`�k�L�������VDX�5��̓~K4W��ZIM7�M�7p�i��o-ſ�����������ځ��ۡs��ς�*�'N�)&�gy T�����E`oM�D�'����Tt�΄[�F?1?#2�C�	��W[?���?�1���̜8G �����(�G͠� ���0!-+�1��>�ȋ�b���r)��b�⸚>���U5'����u)��Z]j�Up��$ʦ�]��P��8Z�kg���Yȱ���l�JP��v��a��|���}툶2+� O C�6��f��]=8=}�8�M��p���ZC���0Ml�#hB]���H���$�?�t��-���˒�P�ںxe����$�����1(��n��(��n�3�����q �׈�X����0�-G�J#�PV$���e/)�s�.	܆�"8OSG�Ͼ�쎃�U��L�m�F���J&=C�6�o�w����ĵTZ�ZȤ2	4���
u[���څ�35^�/���ϸG��f�f��qoڈ��8d���1x���&>]�2r��r[�+�����t�L �j�l鬵�w\_5�V)O���5��_��L�R󖜔!Bt�����80��)��q����[�l;�G;�JX=����
���t��_7���)ҵ�����^���h��EИ������d�XA0�hƁ���m����$:n�3p��L���Ŀ����?����6lR(op��^ �|���K��?��V@� �:�Y�b����6)\@��`ڛ�r|��Ѕ��Q�j�wa��Y]P[�_�qg�ޙ�$�FK�Z<r��3����&Dw{�نwt�	/p<�0�"Ҽ�� �F�1�q&o��!_����zF7�g�~i��D�xI���Rn�0M�b���.�*PHд���3�ɴ����QυK۵�mi;9�F�@���Zu�r%�pFi�1Qp�b�jkU�ĸڅ�6>�*�����#�\��o��Z �����l H|T�w�`����"o��M�#���o����?Se�M<�����+����%�����l���f
).�d�~ً��5�RW%��|�x�N��E;�E���w�t�uQ�[�Y�j��e�������.�#|�X��=N�%�)m<R�ǉ/ȿF<g+H�=��pm��%f8'䐞���k��&�/��3:��ʀ���OS�`���d�W�6��߮/l���qd��8���ؾ��l�üڀ�Y@���v@L4�Bk �Xn�u�����]���g$:�N�M�/d��L&�Vng���Z�SP"������L	��P�K4*H*|�zz�Ҳ�ll�4v�0d0����1�
z�����9�g>0��OY����%�Cм�>�������X��/uC����|ݽ}=�O� 9��9�C���kn�ef�د ND�6�=�yے�It��!�{/�щ��q���lK��� ���uw&��/"�M�- ���,���hh�/����6��l��:r��c�)�^Ȣ������`ZۑY���~��R��Z/�'SDǄ���i�!`��K{�M���������.�Me��f��6���d�x�	2�O��
�v��f�+z�w��&̰T�Bd���1Ю�1S�o[l.8�����]�A����7�>�~���ۜ�}yt�:vu�1�|��Ja�o��\�w/��[ƣ�����%�p�Ԩt����\~h�`�R�F~�I�;e�٦�x���Ŵ(K�����B�;n�@���f��h�d��?�c�r�z�����Y�Pa��,��/�*��i�Z(����)������mXN�U���|��E�si��苶qv�#��o�>tȯ�4�8'�����~~ɡתL���r�8��˦)돵�놜p��\/�ADU�����9<nr�`��������O�'b�b ��>CG�ңL��O�j����)�/����������
�w�bs���d��&����x��:����[}�@���O��޴	SC"�3�N�2s�@��D��ķs��h��4���L��I�τ�MC6�c_q�I�➮�n"l_z�r��"��u��I�:�k3�Z�>�9��	���������D*	 z���h�R��dPGv�`�|I�j,��`�&�cԣ�	y�ng�Үiه�(��gŦ����.�D/��ߠ4T����W$_tlD�=!�c�V�cQ0!>d�Ob�͜G�Y�Y�U|��!P\��Q~�b��Y��8�D��[*l��[�,����VRW�����0,����X�1�×;C�"l�ۦ�
�ɢ��-s��Ǧ���X�@�5)�z�S�pz��E����^V=�̶�q�:,#e�X�����D�Q�'��KwO�Qj�_g�l������)�������n���Z�)�9ɓ�d���#�149b�!��m�̨����L��Lo*����E	&��GL��� ��p��$�9�r�b��dY��JV$����zJ�/��3=q72H�І���y�vZ}�	.EEЕ4�f�M�$*Qx[�C��vD���`{��}7�]���vsw��l"��0����=x�Z�hm��`�45��*��翭Y�t�`JbbbϿV���IW��#�Pml��ϻ���^�\�����g6�x��[��b��7�9�7A}��!n;=�R"wr��e�s�#���o����p��8��Mzd�r2:'8<����S�jTB>���X��ch�4��4r���zx�k�1�9��:7�zj\x�2Lrf��Ӥ��]�X�WwC��<
��	�������)J�L������!L�)�x�1SVzWqZ����3��c��jc$�/� 5�F4[a
5���H�� �{~��7��w�.6\a���4&��,7g�j���դ9;�UC
�:����m-���W5/D|ۆL�� �nm����G����01��|ͭ�Q�sF���E�s?(�ԃ���s�2TC��j�хf�h�������%6d���Ml��+w����$�t�Nd��E)ک�nX˚��o'��>�(�l>!��)Q�^	ڰ�u�X�*�1Z�*�;�S�2��di��5�>��:�M� �)
��O��|c	tflO�o��t��Z�~X�Y��[d���l�^=����`���6PѺBB�#%g�j�@k
o��W�^�i�ߴm~y_f�D����޳oېx�T�!��yf<w�6�.U)�U��"+�-pA�ƿI��
���G[CwS9��<��t#(�x�
ʻ�A�У�k��w �˥��e6�U5��%Y��d���rR��k����+0�����I�Ω=h3R��;9B��P��l�l���`�j�ܦ��#_%�0c�	�IRc<4�N�u��vN�9g�}�
�AڵJ�Jwj`�]n|\�2�Y�t��sҩ�^�v`E8���]�J£��O%�=޾��<m�z�$�Y.�X�6��-Q�����h'`�u[���y�V�=2��F�_d&2�Eq�M?V����؝A����4�V�MAo�u"�XI��/;�= [0���O��VF�44�Y%h-�o���騟�ꐰ���3���
��7�h���s�m���)��Yվ�P4NV����h���{2��`�]4 8g��b{�/YI޳B+�v`���^��}���O�_�遨`4�H��%7�ez����V�ďm �w���<�4H�������c�2��t�?��6��G���c���������7���;��F1�<���@���y��.��Y����,#[�*�4�����-�H��9F���� >�tk���-2���hvu�/�w�|������\,�3��Cҷl�c<S��bjDh�>(�q����.�����x�Q.Ǆl�aY��zf���X��Pj���P���1�υ���n�:ì��L�@ClPj�������T���4�Ǫ����2M5�go�x�FP�P�� ;��L�OHN�O�H�o�Wk���f�ƭ��*�Lf�Zw��ON2�uw	�N_��B�N��~�:!�M�uC�����lZ��T^���f�w[p��U��$���f�~D3o���+K�Z]�;;�BV}_{Z�j%ˌ�#I�`gn$��"?�l7�����?�L���)Z��Vg��k�)�F��ܤgӊ�黱�)vؘ���R�Ҝ����e��Ù ��]��?�ȍ�qm�m����-��W2�7#��ѡ���r���s�l%Ri7�K�#��� ^�^���ޡ;�Qe_=���V�VǗE݉Ag�d��ɸ��
Y�"�[�{1Vʵ9jj�)�?쟴��gO��H?U%]�3�E$�$@���Rk՜�.)�t������-Yr��<��K���oq*�GԺ�+�'�'�c#����XV�h��|���r���+��p�>�߹"lz���~'g�.c��.�b����F����֠���%/��ʊ~eA��zU���*��q������E��ܵ/sf�'�Gs���_j��9w�I�����sKv�K;/{�zniz�?W�����5{�ܭ����o��2�h^Iq6�1�I����K�ȂE&kV���_`�\��}0���ܾZsri��@�����
4�坧uq{v8^�L%z�(#���_��uJW��0��>W���q������0����k)�N{����)H9��]�t
�T6?s]��Y���*[
�e�A��n����Z9x��!��Hc�ճ�g��B�v=�Fe��JC ���_��jl�,z��e܌��%C��{�Q�&�(�߷���(͸=๿�L�w�� U�p�݉�1뷟��u��@��n�������`�>����{�j>/�һ.k3������"3�Y�U���q�B?�}�Ψdz�`'qU�e��fZ�%�9`M�	����9sS �6��() �pI�G4��[�f��.�Iߦ@Q�ԡmy�^�L�IJu��(���E&LV�`A)�O�V�2�_*��O���.�	4J���!K>�Z�3�Ճ u cm�,؎��C����;#��݆���L��ȢN���-��b�j�_f��%�1�Yp�H��H��mc7�nd8ES�v��[�nK��t^,�"Z����0�Y`�f{�Nq�
w�Føb�o+_=��/UW7/y}S��f���-D��s�O�	�t#/t~��`;�&�D��H���G��F��-��a������n_�u��np-z|D�T�3'��\�OPY{l�n<KC���Jw\������2�Sm�7��󵛪Ilԟw��\R�Zm��wkH�d��d�R��5��[a��*~V�[�c�3�1x]Z��U�c"AU�i�M*%��5M	=�#�D� �ˈ�GNi����i�_�	�S�B0��.F�墘�*���路Yȣҫ�N�u�N�����X
�?�R��Ճk�����͂��Cy�'@_����&?{&���(N#���zo����M�0���8c��=n�Lf�|baN+��b��JU$a	$��gz�C0�i!UB�K���4[��B��r�U"�:��?T�����B�]|b`����=��F%�U�+UN�N�/Ta����<��I��q�a�/��p���"���������½
�[g�+�?6��yj��-L�Q��K�0�3�:��"oa2�Ճ6����w�5�˻FiM�P�f3���������xs�u�c����k�B��yE���t��ۭ���/��o_h�YM3q����ޡ.�W-��L�	~˲&�������{(͕f#����T�$D\�Z]�ɻ�-Y"�5&��h4��	��Λ��#2�v*�K�(,OC���:�@����]O��q�z;B4�b�3���䳭�lSD�ҋ�ǚΫ�l8�P�S���_M��5���i�:���<RB�VM$�Nb���P^���!�V�B�'`�d�+`]�_�6/ۉ�F��]'�q�*I`\�L�Ӌ~��n(|0-����~��O|K���دCb]��5;S����.�����T��}���=��k⌟�&
t��he�kJ$e��d�5���[ә~g~ ���)cc��������񵗥�6���زO<�T���g�='�]�@����
��מ	��-k9'�fh���F�uT�a�/#�. ���Vݧ���/e�{��(>|����	�vZ(�����9��X-^�i=U��i��~U�`������W�|[�=y�ڲ�A$GS�b��MpV5~7K�T�&A_��V "v��[�m7̭e����C�����ԥB3�i�c81��uժ�`�
�!"��ͮ%k��[��,�fR�)oJ٘�_�����v�qd��=�.Rz}	�rU�*]L��,��'P�>K�M������Y��7�'_�&{��X�"+<��O:y���ß����&���Oj�<�k�s`xz-1���#'	S��~�J>�<kT�o{��3wnV�|�#��C����?V-p��ޅ��N8�����1��D&�}�ʈ,�{�h퉏n�7�0��� �� �Q0���Hc���v�V��	�7�^���0z�JwF{(�:���iOi1��K��+S"v���Fܠ��<A��~Չ���	�)�UL��5[���:�M�r���<?vvrrBU�$���_����Fe<���V�0��3T$��<��#%&�!����P\8-��{��7A�X���%�%�!o`��5�6`�}����j��ѧ��?������V��k%XY�^2�̈́�/6�f�u��~��/��IəZd\|��B��>z_�^�(({y2�4�)���赀�^�-O4�� |A���sb�ڡm6����nZ�����a�w�6���F��,��?�(�FW �� H�sW�D+���@M��ք��O�=��@�$%j���~��0L�������oM�A^S����`{�����p�C�a8S�E�jH��B���Oh���Bf)ڲ�v�7�Iq�ឍ�]t��g�f���1k�5(���kr�����h��ճ�sQR�-�"$�`�к�L�w#}�AC��K�Y���QOQ߷�@�5��}��j�H��s1N"!��D_!s�����W�D�
���P�T&��4O���J����w�&��B#v��h[�KjބU����\��[$�)��Y�c�kP*<��[^�IBڇÊ�W���G]��$G/N��9����=�G�;�)* ��B���@}t��]ik�X-(}����EE�w��Z�f0�V"�!wj�k�1�t}�悀��Ÿp��܁�ˈ�~�����_�(5[��E��M�j��U��0Q���@%Xhm)ve�n)���Į_��H��v�1��?*~��F������DJ���`��M5���������IkZ�RG7�l6o�͛w��gjs��:�8�%$B�z>AOǅx?�y�F5�t����b�O�(G�v��n��P��D�j�����ݣ�l1gOC�c$���uWI_�}�����(̣�Z�Mʛ��5&�� c�O6���E�s������tf���7��޼��,�qq�:>���vV�4�u!
ȓq����4u4�c@t�)�Y��w6g�3�������t�"�:8o�W����R*j�s�t���}��.���Gw�5�{�pjy�I�;w	
u�k�mH����c���"�CNOb"ob�����2d���	�� !6��4�32G�R�S4MSk���� D�Zu��s�گǋՓz��_#>6��]�Dbp>M�*?�ߨ���Z��o��@�Q��Rw�C���1Xt��}�
]Q`Ndi�@�����Xw��yf�/��٠t������W?�R�Dq/�o�G�O��:��)��ʮZ@�9��y7F���Q�Fz�z޴�O0&�G�^��]�}�Z@U����R���H��+l�������aNo��_�X���`B�������a�p5s�:�ɖ�R8����N��/�sw�uTu}���(`zy�hA�rE2ǔ,M
.�6�'���&@ �/���Uœ�TTT���M���B,l`/�moHm�Z�ߦ��K}5���wO�ݹ�u�A�v/,�)�8�_[.�'�NE{[fP�>�J(�n�(x�Z�,�U۴��զ�}Ս���éU)<y2mA��
�[�v�a�����B\5��g�2��'am�-j2UQr��V {���oH�{�"�!��J�a��(�V3�!E��lm1ºmKO�![
Z
O�<(	��M��I;޺�vj��5������w�?�ە���Y����o��0�����m��-�c�������:\����T;z�?FH�i ��-p�5�C�3	�c���a�<���*v[��2�I���
�ڎioɾT~��p ��pv[�a0|�G�?l<������\�ɀd��tA���h�aP���Ξ�/��SNci��z|_�r��f�ٷ��4�尧��!�y��w=�y������`�#���!9�kqĂl'���#�����RJ�ߎ�ɋ���>��l���jg���%���̏�W{&���~���ygښZ�l�J�n�n�5��.+�m���dYj�`q�[�N���=��K@[J�k��L��Fl�*��Z<�r@�o�}�)${´�a�k�p	YtV����[�(�dq�y�������[H?#�\-lu$�K)�
H��W>�d�")���Y��	�R"�
��x���膶A1�0G@����.)}~Q,��Mx�9�������{�z���{�����L��?�^\�`��U�'"�9��ߵ���E�zP�gԀ�i�v�!���"MM�&5N����W���f2"��S�6��`�5d2��?�:�I��Q�<�d��܁�qx���G��U
w�Ȝ���k[;ƴ�$����.ѻi!�_lnɩZ���L���mzh̗
�N�J1�D�'�Ϙ8�����~	�a�(�5���X"مs�Z��/n߭�V��~8����)�W��B�\��d�$r��Tq6U�I�޻h��'e@O__H$�h�˛1�	"Q�4�ƚ"������ń�^1��]zXIQe��i�'��/X]������t2��nr��^��Ǘ30��P8���/K�2�D=�T<��܌8e�c3�k��;-H��C�rS8��{ǉG�z���U�g�;����8��8���>˰R���5���������������[�-^[���IM��6h	�����y���!t�I.�����G/�;ϥ��0<�?gpQª��Ղ��N �J�����+�� ��68��p��;z�Ɩ���W�S����0ߎ��~���_�����cev[����[${ ��>i$�Y��u8���)ώ�c>rmd/#�sK�B��%%�+�nt��d�H��ӓ0ni���
¹���uM�I��~��wnj����ou+�o.Z�eO�uf/S��K[iV��z���1�A�<�M	�ǷZ8��j?f4�^W� _�\���Y��a"v��錎�v*|��i�Jޮ�	�[��6�'��[)~c���_e׭*1L��b�/Z�U�fد4�A�!-��h3e����J~��ث�b���������?�O����d~�J�mL���s����x/u���i7q�~�����.R����2	���I´�J��9���fN��U�������t5��Cl��}*M�����F��'O-���U�x����>_���O�qrB����mᣠ���^onY���|�L�C���W �����+p�3���c��^U���I!g�����}�l��L�?��4[��x�����&�f�-����m��(k�a�Z�R����/?�3�\��vi���)���̶ 7Fkx�D�/�:_X���:��k�����,im���z�C�
�x�P�#��-��|˳g>R�`M�&�L�������l�F�߶��+n����(��3[�N7l�]-���j@��{4��%����6[��I��s��'�a����}��#zp�A-(u���c��Ǟ'��y}ƺ�fPm)�Ws��1�F��z'�ɟ�x��u��ڟ��Ơu~����+
}r���b��m�z���}�Ů.ݍ�`hT��E��	�,�Ii�M�����-��m���2��K���o4PF�w���Z0q�������{>���l��B�E�(y�v	��GE<d'1�tК��+�w���B�y�Z�ϣ���΀H�����ѫ�T��b ��,ϮH�4C��Ee�<>�νL�r�7�?�p9Ļ��z�(`���I�\����qgx�]�+Nf����2�u�^`˙W޳ф�C?6�JƦ�j�'�����=�d�Xh���B�,B�H9%�)M��]�r�H�d0�6�_dv�����ϟL��m�a�3�KcD�w�)R�x���\w����_K�ڈqhm3s��hQ��߇R�(V�p�9EgZ[��μ�#o.?��WO]�����a��S��Z9��XsQ�#My	Y��t@UOZ��W;�3��Ub�Q�1�L�۩X�#�C����a�hZ����Je�!�+�D	�;m���C���ug�w.�F\w��H���kd�KǛ�N ���(f��z ��C����@%��D���u�z�|l#�<cGS�?;U�RP�Z�賃�{
��|�����I �����)�ˌ�ي}\�/d]P+	��:�H��a��OG�W��r��A�ese|w�糲����n�׍^���w �~4�WSW�bt�	���aܕP�1����tw!	�å�x%���?fIM�e��n��ƦAu'}ME|�(װ��4G7�H��TM����W�eh66=��0�o�1�Ю���-�FBD��i����"���w�ќ�C?��(ȗ��^��)L��\�li�I䢱����=�%�W�dd�lF�q�j"�W�(����Q����I���쿹���r��`��V(��9L!�
� �f�m��5S`���L�%$�T1��6=׿0Q�lm̐?�5Ef����E�MY�~�G�hN.����k���>aJ*�Γw�����1���0�/X�h���{�U��Uu��^�����%���T9���n��'���2�D���s.u9�O"��ʸ��#��+�^��=G�'8��&�@$K�AO:�R�"^կj(� h��`�/�ۭ�^��hi���U��q��D��߄O;Y�u?��z�g&�,�S��{qJ&兗	�Gg
�쥠i���F��&��5UD�C�!�#R����������T����ć�!���c�uy�\���)�Gx���:��W�kP �<!���$�����B��&�9=E�q��2^���T]`%#��Kf��	�Җ�F�d5��۷���xe��������\��z�o�\s�'��[�(�*�:���p���@
�y��K��� �1�
Wvz���XR�a�OpQO��{��w{	L�̀�؇Ď_�J��ϟ��9��p4���|	)p1�Ic4�E����1���攢����m�J�Yo�gH~���Ʌ��	�Y�9.�cs��?E���|K��9��iZP;�f��������:J@�B�U����������H�veX��j��nط٤[\�R@՞�G+>�`vIzO���� =��pp.��R���Ԥp���zSt"���3��!�KB�.X}��sQ�d�&wϹ�M�1U�i���#'�Q@�_Si��t�4u���|�ΜYh���
p~[��K��Q��*�\4��c�R0]��L�]=���ݩy��.壁�Aذdw��v\JCI�}���	��"�e���A��e��l��K���@�"vƜ�����UB��e}.~S�$�Q�-���ͷ��r����2�2�P�k|�Z�z�M�O��"/@��r���v��(�]Ϯ����f� ���C��Z���@��>+���^g\[���A^��6�u�[Ac�� Βc��}G����P{L
YFٞ������si��� y�ú�΋�_Ek~���kaS"д"K)_�tٙ�ʼ�
��ݾoF�)V���ӣi}��"l I�9����a%8Tr"sw�ߚw8����\q}?\S�l�zL�ܸ
��k�6�[�����í(�� �%�^��>n	!��Ied��&X�>β�_�m�Y��r���zB!��ػ��,����J����IWt�F�1���4��`�u� �@��K�r)82��/:+
���,��g-k﵃��	���E�O;N~�ߦ㍢Z��C��P�bݘpI���T�j�l��-��](pr�]*�lU�h4
��6��GdtG*Ċ�Ԙ�a�mC	]W�@,cm�,S��э�w�lJ���ܫz|�TZ�{׾�X]���<,�2���B�s�2����Z�%��n��R�����o��)պh���(��њT=��s�z��[=���:j����>~~��<��~���ȝt�6�B*-����y�m������
w�@�!��#?w�{��?,o����;g�^���B}�G��b��B�e�"���6�d�n$�yj�QV���G���x�<2#���A��_�ܼ-�LL�ON`���Gtf��.�u䨹��Z��E���҃w��%��0��g:���ԡ�#�]�1�B��6��?����	��@x��D��0*j�~R�/��Ĭ4�:7r0�v~�И��f`
�n�$D,��%2���c�9�9�$��9p�RՋ=R�����q�/,}ƕ��Mwެ��Ђ|X0ϒ
�Qͨ��Z���UTxc�.�a�z�	���K������t$쿝#�K9����I�O/���J_No!��Z����B��[��E�Z ��h��^_��o̮��X���y�q����ιݧ�#���5���:�W����8������o�4�����F�.@�V׆=�o{'�TE�y�����y�t˶k���;)U� |��(�b�&��3���?��>�\��tQ�K�D�Jr_0|r2�Go9D��)�A�=�:����5I����_(�`m��ϳ����H��=��º�=�<��m�"��R�:�-�������yF��b�51a��4a��
�N�i��X��.�}�餥A�n��I���P�g�X']�.��;�#�Sk]���`+��*c�[���-�.\\�T�&ި���l����|z/�Vh`M�
���m�0��&)�~d���ڴX�Tr��Z;���,vw����M{��&�.�-�s���������5K��g��(�ߴ㊵��?��?D}�C�_���HwH��ҍ���Hw���%HK#0Bi�Q@@j����#~��}���ٹ��Ͻ����1�Qw*qV��T�WB����Gp��?S�6�hb,͝���.��[����}�Ƣ;�y�D��ey[K}��3^���Ӛxk�F�no�:�l��H�2]���������Z�{�����B���U�1u�ƅo� ��AQy=ܪ�
�;R��~�a���RtR�磳ŏ�:��A�h��â`+����ǻ��y(�Z��V��78?5��65�����[��8"4���%���9{�+c�h����~�����㪽Z�P���kV�h��46Ƶ$�Q�[�j��!L6빥jo��J�`7���*��'���������_�.�u_�}���gF�^�ٯ=[�K+g�!�I���R,;����ߣ�QJA�iU�J�
߃7ݛ:��1�n��	���f0�@4<��DW��X���,�i�F9���q/y��C�P�o	�d��&���
�b
��w~�ox:2~� 9����4�ڮ�Nת6�
�nJ�NdI�X�m��w=�˳���ݞ)7ܫiZg��2�>`ˇS�T�n�jl�J��n��#uQ`��T�k��&
t�=n���x+�!�iį��%���}�F�q�V��8��45�ڪѾئ���Q*(������_�9�Ȳ�7Q�!`�>0���a����r����WM�_#[�b���]w�͏mz�%�[x 4ި}��ǉ���k�A����Y�Xf=���S)��Y��~קPC���ˏ�N(�Oa|�r���_���GK[��+�au�jc�PN6��ܱ[�y�ޅ	�j�� ℏ>t���C��]��j�4�v��xo�T�B��=Z
6�J��)���Y��E
\p��P�V�����Afg��m�>[�$�9̓e�F��i]�2D ��m��S�S��ˏ ��-����,�Qn��|�}]��<w��p�#��U+~8QlY���*�?�h�o6�V?o�6Ҧ�a/�>�ϠA܀���+�D*�7oE�u�ju�y薿+�奛�8����e����G�#� ����^&�B�]9�R��A�o�מ%���G���j1��"@��o������.��F�΄A���~k6���1j' ��bK�ܕ���~���.��'���H��}J9��<�\�yw�J�Da�V��(�J��O���^J���*rfQ���x����D��D&1j�Q}���Z��iSK�'X͉���9A+�����-$AĵU����ϥq������<0�!�B���_�IKzp�Yj|ZMhNt�����-��v��1��f9�/�������O�F͸�dS�K�)&��d+N�b�J�G�b	�;�#��z�}_&X�l6�7~T+N��ia/x1�bлV�ld���v�]Q����x�BO�O�C��̑} �nB�;��뒞�t�ن��X��/����x�+����w���9%W�Iq�M�Ո��9pU���?b��ʷ��j������f���6H�X,[^C~9�j� �$Z�G^�����̼���EaW��Ȥ�+Q�:(	q������4��Xqv�}q$��m�ɣ���?�ܞ}~j����ϼ>��G�+Y���c��%�Y,�R]�L����*�d|$̬AO\�Ig>[H�6�hS���'WԌS��7F����}�|�E��Y�B��4���w"�H�L�r��e>�7�#h$��)���\�5Gl�c\�>w�,�F����KݗT7g����������?o��Z�ϴ޽���`TιR(���Hz��f3��� }}xݸ�>\�9�&P�U*��=V�S�xk^j��{.���!�@ۅ �O;			�n�W�>�&����
��ݭ`�d]	�L&l�����,��YZ�S����}������"�8�%�m��Q�D6V�z5m��vJ ���s�V)/Q�J�l�\0|W�MF�[)I<�����ّ8�o���OO�GĂߢ�m轷h3�x�_��%ާ�OYG���,Yxq��qJ���7�?�(���U��u<�e1��}�2����"k�]it�~�#h��'��x��tq!���/�K)��`����/��`WbA7��;I��=7�����h�� ����z�ېo��#|	1�C��o�b#R��|:�#�hM׷�S�K�X}<Ԇ�&.��4ӯyEog�M,a���[r�[�<��7�� �@�:�6�v]'iw���:��G�� �3p������]��j�Vm�ʻ�°9G��j�h���&ǚ��
!S��]���"ǎ����%p��W��_�d��!30����LB�n*�b����~��T���8r=�K���腀��x&e`�`Ni;߷v7�"i��v�	����U�Քi�7�y����1Ą<��|2G�+f2�ކz{������J�#M��^�6f�c�$�l�?��z�@�
���\��,GUb���Y�:E�����/LsD���Z2Q�/��bz�t�(�{�O���"O̶�>��|�f��;�����Q��\����T!gՎ�}s����4����V�'�y��a+�;���ʚ�g)���ge�X�H�zԠ��L��ˣY��7���L�]�;P��ޡ�9b*u)�9Z��%8��dLx=&�p9�x�+
��>m|a4Я����#-[vD�]+C�E�1�*V �%,��,
c!mm�N^LZ�kA�k��/6 �EE��Nڔ8һM�ǔ=� �%с�iv���҂;mQ	j�D����c/ϭ_U+>�}߶��^^���t���!�82?pw���[#�x�z�m�x<R�%wM[r��c>n���ͽU���[�9a�͝�ư��O�f��3�U�M�ir_?�MM!�����y����j����N��
�;|���%7?{N�E����Á�>h�v�tǺ������#�Y�� ,T���ɏS6�����`&�#x�ɒ�X�<D0��Hp,�3�sٶ'ku
���R���#�#�a���f�7���B����$���񫳰����F�8����q�{!�%���7��}��hDa���@ -A��Z����l��9d̟��n.�
ɷ���{��6Pu!����fh�dp[��f����޿q����s�"������� G!򻶙<�~��������2~=,�a�=!�k���?�|�B9 &�D���0�:������`�OF��'Е�H�þ��E�f�@�,b"�ύ�<8��Z���X^�J).Ր��M9���#��u�)���,�>��2����ɼWÄ䩂���b�3E4����y���b���n�tW��[��wx{N�4�q(86�X�%�f��#8|ʶ�&-� >�߫�%
��٪��Wj��4>�7L57^�.��-
� ���?��Q5��	d����4��v���$3�f�c@�_���24W"Ƅ��!Cw{���w������� Zt-y+^`L�+Ǽ�bɔ''��o��ױM��1U�͆,�-��\���v�Ǿ.:�jN�)ܜ�'g���έ�5���1@�9Ύ&��]�5����{�-���&�R�f��\�%�ꓩ�4���e@Ց���4�ܗ03r�.hp^��e���筣�[����!�(T��m��P�=i�EN���u4�$$�ǫ��p|��/�%�A��rv�n�������<�1K�?冹�ڊ�&��̚֎16Y����6*]ND#�^=� �2��Q3��v���cvӓ+8�Pg7{X��4�L��Ī�_���66�aݮ���K������Z�
�J�������3��S��C�GP.
����r�!��X>�骴��Eܰ��(���.m_I��\�W?�����MP���hc׭#�z[%��fDbO�~r�BAf��; �m�}���% ��7��m��TOL�*�+���t-o�o�;�
�Y2?��[�%��&uX����׾���~�YܘY�߹�մ�n�>R)q�=�����;�<!����]K�f���`�,?�����42٦�|��R�.�@�z�-�T����H37D�}�%����2����{�������5˂���f!r�����XU#��W��6��+�yH�gݳf�-�1/����9�g�_��-�Uඛ�D�;��ň.V�n�C1�oM�T>��|��o�<#V
�v��l��S����k0��K˒��n�T������rAx}��>"|��~1���^/�?<���L֫��Cͷ0P�{�ogQ�Q(D�όpe%������^���"3�#�S�^M�y��cnc���T=}l/@h̜Ou���L�$uϭ��1����:7Aˇ~�vLJ2�$Y"b\ԇNѳ��2����u^� �5y�.��`��H��F��(�`��l���6g��C(��fM3$Ǆ6�
1�+�wG_C�
�wA��.���8@=�(��� �÷�wUp�� ����i�s<X2#\0Ӻ]��8���W���6�-V`7!�i��v6��8�9y!�u�R�!\�g���#��&�/�NXӚ%��&��{�-�~��	��t���A4hgB��Q\)���c��!2N�N&� ��6�z�̩�Q\��F5�Z-�(ˠ��O�[�9�<��7K���r�7;�g�ΏDH�=3\�g���w���iIm�Y&�yq�^��\�������G���'����	�v�?(��F9m��F��>�}U�7O���(5�$(�gN�/��/_�֭���_3��<9�	1�kS��z1�>��6?%pz��]�B��ԷY��������h��Kp}�E*\���,%��رT�J��<���RI����4���P�L��a�>bŠ����8z �j[+�.|:e8+��o���ɴ��#���Uo!�g'-�bPy�g�^�w�<9?`�O��Dzh�4����J�l*��̦u��(�����M�%@C9i8
��Z2�u���{nI%���!۴W�0�yB���#Sґ�O�al��f�~�4H���H4�JP�����
CL�R<��1"�����V�3B�Ww�h=n�L`��8Wd��!�v~_��vJX+��e�� }d���Po�b����t��� '8��[�<��`��»ک�r08gAUHٻ�$�ܒQ�����u�c�9'�@�G�����M9{}m�.�WO-ѻ�V0Z�2瘘֐+)��L+ˎ�%l����yn�<�eXuuuEŸ��@���jV��ɠ�S�z���!�]z�E�2ס����%9�\��q�48�I��c�T�,�]�{�^̍���j�$>��T��t��/Tǃ�Q�D6�v�u>��h����h�._��.�oў�i%Ɖ��i&�B���w�v=��'��w�w���%�����Q�{
�M����g�݅�n�H�[�B�dw�ƾ��w]rfy����uகX��/B�W�7|���ܜ��;I�(�H�D��+�Τ��{N�&V������!�D���{�U��)��0T�b�W���(j���S�����8n.�.����Dp]����G�zM��5���Ds�mj�;�B-����s�嚠���b��A������̄KY-l,�·o�u
�����t:}���ת�W����T��~��,�>3��)�'�i�F���0fr�3���4k��4��ڵ1��<�,��Dr�1�v+�����N�;'sp��Y9�������œ��5�M(ߦ����Kt�i����n���3��W�.��su�e1�}��xh��j�����&x�~���-@���-�V)��L~�'+�4F��sę������}��qp�����VV�F���p�i�hO,DK#�Q"��>jQ���d�좓�E��C��l�j�0�-�o�e�r��Z�m��L��3rW"���q�kB	�G�1�%�%!��J,���<���g��l��<נ�B��A!�m���*Y��!|��̄������d�΍�M�:�Ĉ.>��B�n�v�+@�9��5�e��i_q$��>3v��C��l���������Nѝx-^O�&y�Me�������������Z�)�����Z.�g��2kb1���-���>�6�:�|��V�������W�ir���Se�������:��+Q���ȟ�;<����|{��g�e�嬹�%����7Rc5~mf%y$�xL��y���>�\/���<hjQ?��#`��}��p�>}��W��K蟄3��V��ޠP���"-��њ��C�ʾ硸���o3ǡlC�<�}Gg�cTϘ�l3�S�o�3��yvWbփ�������������W�
;�Ǟ�A����U����y�?`�7ʛ�8��c�J��錏���g+I0��}��[e���<�#�M���1Ο������,����t'��������qu�6�/�Aw�,�� ���>5<�f�� b����i9*��x�<2ʆ�\��N����B:��mx =�G ��%	"|}%C�7K�hޝ~�}�N�,(]��9.��C|�{#I
��b !��t���Õ���`��iB���p�����h`�,��w���K˒J�ar���7O�cnV0�ͪ�ի`�b�o����^c�#O?�S>�4�.�ߗF ���`�-KJ�	Y�i���]?s~>)�
�&�~���1�(�+�8n�x&�f4��)5a���6J�*�r-g?�b��	��nk��|����?��-yZ��LGi�(��>�}Pڽ��@PR�[����Ä4���e�z��;nYA_裷�#@�u^�/�',7B9
�T��A�}�S)sV��\x�6\�o��{u����ڵ�����]�H���o��Y�4�a�p��
���C�����g~ۇ��xt��u�ѬG�)k�	Θ�v]�zQ��8~���:���Vk(�S���q`���u��.���7IO����5���"��ݸ�i ����bK��#�\��D$�h�uz��>i���9jmo�Ӑ��3�C�C Va�Gɡ�c)�X,'l�_9���`���W$j��VŉK�:	�a>@1W?�y�+8�KY�^���tb�1�{�ڒ�;�n%�W�����j�l�n.�gۣ����˷s��tu�* ��>}R�kx3�0��U�Z�<]�&��y���j�-�R��"k[Y7��4����l6������q�B�'��3N����� ;�WCq,���ߡx�?��k����]�X���t��?9vq��\e��19����AB���?J'ۡ���n��U]���'��rK���B,�-+ZO�%Y;��A>����SM8�����o@�`��>u>z������-nP?��4:T���#-����,��d�J7���>�k�4�u�0$�=D#`y\�5\�V,x&1������5��Y\������0߼E�װ;<���R?�b�#z�/K�,�t�z8�'gNB�l��;�3)���5m|vfq�D�����YI�]"Kw�����Uɲ���qB|6�8rL�X�H%�|�������a�kn��yםe���;��5aj��~l��b+Xʵ�c*<8��=B��/��;���29`���[y����U�B�\�
�wF��N��w�Қ�n�Ar����J�A�:&83Zc�i����:�9���9!g���"<h=�>i�����_�V[uZ��Ja�PzctP��#Cu����>�vq�+K�}����.9��}'r���c�.�ߞ;v,��ڹ4,=n�����εa������qd��h�r�\Ġ�����`N[WW�O�?��w]��__J�X�
�elX����[ *�>�P�Z�	�$�׷z�̫ߣ���s백=K��(I.��cET�۾�7�?��Rj�T��g�m
Z�B\�ۣ�-db���p�߽~�6(�i��ҽ\�~�Ot��B��b Q\�A�ū^���]妒��>�WJVoS%:j� ��T�8p�x��a:g�)<p�啚,��©�CA��E����;3Ä���F-LM������=Q��ח~���ah�_L��)��u�,ٻ�w7����]�S�#�P���}φG�/��ϖ�/|�0��8�E���3�����vm�=1,��&7��ˇ���ȼ�{��q�����r�/ͮ+i�7�����&U6�cy>��M��wK����Ĳ�;~��%*u}��_3�����V�Ƚy^���FH��j�u�S� a|�掐�}��@_����y���l�ۦ1�jL`�v�s����4�2��6,C
��g,���C];��YS"��C+�qe9Ø(pR��%������O�Qӓ�%��-�x.Ó', ��]�Ӂ��7�˲~!C=�8W������!�SZW��"�|�/O��6�J�	 3<�C75Օ*�|K����6�[1[�l���C��tg���2��o�0���Y�:HuE�[R�;qoKp���R*��Y�����_�������[���C���]�YB. 6�_
n�tB�2�;�j*���H$�~�� ���<���5Gl���^�|�})1�͡*-�{`�v�S(D��v��9���y�a�) {fKt���NC�~뎝`t�uЍ#$���L,�;'� }��ٮ�{8r!Iu�dNq6
ܬ��)����Xܹ��C�ֺ���Yϐ�����c�?�'�Z[ˏ���߈�/��-�������6�^ط��	��M7?B���_��pgD�|�W V�\�V�đnX�pN�{����-����B�h��_t��g
?�n��Y�����_C,J��	���/�T�߮~�^X���/��S�ׂN����Y�x�<d���^^������鐫/M����/X�M�P.�=KL}��xu��a���la�Q�d}��i6&pٵq��7���?a~��㧷2���GR;7��f��>��'r���2.b=�UC<,�o�}��4��H�M��*�� �:��p���Ql��S��o�0	,��?��-)�Q��/{���9tv��D��4�P�|�0�{�rʧИ�#�O5u�˫�K�(t�8$�E�x�W�Y[/�Wm 8=��w�۱ b�R��!~�iV�<}V(щG&����!���I�Z�@/D�3M}��v��x�� ����
����]
���$�K���Ds/
g���US�~q�cOK��d�����QD�Í�D�k+[�3�R�Co(*l�t��]E7�@���g��%�'�f⮄caƇ�Z�+e�F6<g�Q�~?�(���o��\����憐$�\��ƌ*YO�g��8;�g�/}�@π@d�ߴ�i�)�:�g���!'>٬��=\��������2{̅:�;�,�<uZz�k�@���,yo+�a>�Z��0P>�h�8V�iI|�e�Vi���_��ϖ:�Y��Y�H.�>h<T>���ؗX��1 a�5��;V������]��D�B��ls��v7`���:�i�} ��p�{ܐР���u�J����x�����?u=�s�E͡�/�T�S<���7��^�7�9�!j�9�%�9���k%$�0I.y�3���ս׸���V��~��A��"�Y��sC�8qୢ�Nn��"	��l��0t��cV0�ur��6���m]	��
��p{`=`�X������?y`�<�K���^���tPx,l�/�&1�z�ǥ]~���X��^�|uv]��H�L�>t��r ��t͜����|��7��5��?����t����b�vJ���~��� ���z�"w�{����~$������0���ZY�»�8������*�x�ު�sd���_�s��(z���:N���L~��y��BYq��P���@ŁΓ�_�l�3�El.'�����{dԾL��:�W�"[�qZԕM��E��!�4�T���Q���yȕ_��3z!:,X�B���\x.SZ>�>�"��������r���X�>��
�NI�(�_4+��7���h�1�����M�`#օ����mc�X<����ٲP���1.{_+���|�JQt�[U�t���~��X��V�3��e�ud&Bǁ�L��0u�*��K��l9f�GKM���^cB���P/�>���N����A�s�X�]�Ma~�Qƅx{�^[;'ٗX<�yӾ�[����N�"�/K��4�	l?��J/�i�MЍi8�6��!�kq���x}��aX8���9��O�}��R��*P%�̤�����Ӂú"J[^I`�`*�����sD�M΁Zk�销dM�)��p):�
��.��@d��ϒTӔ���[�0l���u���)(��� OuS�5�d ���3��ІS��A
9�*�j^'G2	�t����4��ZeO7H��&����'^�E<;�����)�I'М�����=^�[x{��6��؁U^~~ϕ`7�s�[(�A�K���q��&� �u��c��#V���"���	�{�t0g�J�=R(�P��k�2O3�O}�M�d����]�#���Ɖ�/��r�1f�1�������ފ?��~�{�7��n��i/��ÿ�d=��"!)���V���?�I���j2�hB� ~u��YwG,*���A@��ר�V�5�0�P��_�΀�yT�,����I2\P�*�+�����T5��Y�uk2c�Hm�5D�ѝDL��u�
���-���
D��a��o��x!��Y%oK�a�6&c��~�{q�;���^O6�Հ[��(��y���Y��+�"]��36��p-������Q>��B6�H�\&f�8�t��Q��T���"77T�k񆾚��{�4��P�Z{����r���(G���Cj��2M��G�"D���Ͻ2{��;Z��R����Ƶ	&:��w�?أK�àa�8o&m����W�ZC�-���$+o��zT;M(T�2��!�����K�ӱ�Y��6�rڒeD���5���#ڪ��YU�h�e��~r�d��nQ}��^�?�u�d7��au�S̘��8�:��c��J�Vi��f(����΁�ņ!Q��Q&��B���?S�F��(��W�m�I���3Vp�oz�1�y�� �/^�]c
�
k�ϖ�f٣��~���٤�80R�?��]�&�4��ـ�j�Qb�@l	KǞ�r��K�Y��>�^�I�O솸�W�y�>(��ـf�%�r����V�+�3#�5��������%� 	��m<�YO<;���?�j��u��uP8�)��ږ�%�'�x2x���|N��(�l5�X�`�����7�yϣ���c�-ڨ��3��D
��{��c��q8a�6�ÔL1gR�䕊;7ߺm$��>�if����թO�������ԥ�"�.��Z�W"dl��	���e��3�Tt�:*�EC����m��u��\��ڣoBb�i݁��Th��&����q��/e����WP�{SryKBmۻi�&�"0�����xk�E�[x�z�ۈa��K�d�`�h:R���xv�B|�^^N2I���C[��X�߂W�(�ؼ���WI|���]�
ݾ�'��͐�N\z+Ι�Դ��X�x���� ��}c�񣆹�68{�jGF����F�*�yΣwg�I:�=FX� d◡|nH"�<�5��{3��R�>���E��4�T�v��+r�=F��ADσ��jR����OMU���:q��eҡAo!?]��<m�����G��W��آX��<YhD�G@+54�J�eL�%��,��-�Ӓ�*nֹ�TO��Z}���&���˿��E��p�r�����x�vZbY��
�
5�"���j��8���`����m��Z��F匆B��=����W�|@M�܎:�ÈO΁^Cee�ɗ��P��_�Q�nO}�bD� (t�A��ǘ0?��'{f	�&���Y8�i|��~�ʍ�H�y���)�W'�$�v���L�5�v�Ԛz��ć�K	Z���1��*n����iNX�D���}��ϞO�O5�
9��yզ�a��Z�����.�|S/v���Y Lv��t��+Z�>�������V�@ ��7.�%�!���-���|c��G8J��H�_��@��n����\����]�j�KS���=�	8"3���\r6�Z
|pcR۵���S�C�y힪�g(04��=�d}�=S->+���ͬn����~���{G���V1\5|7�O�i��!�\5�.!|rRGBJ�٥M4�I[Z�.X���M�p(��i����c��;|K���������Q!;�j�z�����pZ��X��x58�+�6+90x��r��t�&>����m����r���+�G�\����f~M�hw��/�N��,�,��w��D�Hz~�>�7��&�?+���0Mװ�a(�pS��+�ey}|CU�qI�km6gV���j�S��*����WP��hA��
�3�����e�g:&�g�@�ڃ��n�K뮖�,�8��*2�[>��$q�h#cr���\V�Nĳ��~���g���f���'Jϱu��M_��#�Wy=���v�Yy>���pɺ�S���.ol8tS�v���>��ES6ì�>f���`! J���<���y>���X ,��:�󕵜��Ǟi!��Ĩ*l�v:���q�,4!�/�i%��� 8�ִ5�I�>������'��d��=\�u��7pm�#*����k�n�$>Ko��!bԮ�f!���/C��j�*��-؇�@��H��N���]����GO�Og!N/���@���ֲg\�� k�a���H�:	��1y��k��e����g�c=��~��P��T�N�r����F���dE�n���dH�<�2���I�]��h�Ǫ�O�*�{/ķ��H�P�#>լl���[��䒄f��)A�Y�۬l��P����x�-1'�/]0�#�sT3nn=x��4�ͻ��L�f�t���W:�p�h���d镕�w��.�v����)�r̰_!����ׂ����nEWx_ߴ��PN����3���֐�����Sb�|@�x��W_��خ�'�j�䬵6��b�3��f��M\�-H�:�l��y��T9F�CH>L���p��w���> ������*:JK�*�n%��z�)�е���j9�s+0,��=SxZ5�S�����/�9qC���uH�=\$vY��΂�>j��AyP����Q����":��GxN��ŭ��5���3�I�i,g�\�ܻ�ar�&Y]���K�	��"�D�\rOs�ʵ?dIv-�X�cE<j�)x(�������!{�N��L���]`�1za��/��r�>s�`l�3��oU��R��Ѵ��~]�l�Y�緭��#d�9�M��.+�������.��J221�~�!�}ע�&�|�|^V��O�f�\+�ajQ� ���"��ߴ�d���W��j�����>�w_��a0ݧw�g5(۲���gO"w��/���~䳚\�Pf������'��F��*j�H��y�q������c0'
�m��rUw�8��M.��Ly�+��.[]�t�0o��6:�\�,ND����ij�˦�K���g]����.$uQ��?"�c&�mD�"���/�D���ơ���q�r1��m�4�����[B(���o�^���MS6��0)��am"��N*V�.A�9�'&��yO�5�&g�o� �����C���R��k���}e�\�"п����15%��,�r}#�(W�u:�o���6�H4$"�����Qp��'qS��8U��,�y�˹�q�t߉[[3�9#�I�Ͻ~,�(&��^1���ӡ"�%��+����%�Bl�6�|�v��`�@�@����7f�6P���c2��V�d
ѓ}�����A(m�&��c�4)�nN�Y��.ͺ85�{AQ������INn�,��B [^�c������VLYc��"�s�κ���s��2����I@d��}3�L1�"#���^��C���6��⑋��ㆄ�2`��9M��;�`-�Ǚ?	��+��3�ڎ�W��7�\\z�<�Ӹ�����&U/�����{	nå�ӊ5K�o��U�Eh������%`��\	�Uǔg'��|A�� 9A\u�%��x�J��s=o�(��ks<��;�O��!9\S��!L(}�C�����
0�\r܃H�������Y��:,IP��9�P]"9��+��M�ц n8v!�1�C\��pi���V��U� tv�k] B�
1�`�n��,�ۇE�����0B�v+-]J�s[�.�ej����i�3�IL:�dkh0:� �:��<��D������4�L��Ǒ����D��@���X[��*6��W'"8���Z?Z[?�R���4� ,��y\;�G̓D���XcTk��K�|y�ګǳ$/m��N�Κ�޷FL�!
�H�������#M���ew��E��
�Z��t[K�G���s��-ē#�ڀ��d�	(���7���-A{ySb&�ۥR�י��/	~hwuer����8^'WZ�A�9f�����V�9�@ d��O��8�	zT���^����9P�S����h�s,^n��>��F=��
��Z��j��2\=oY��wc)���;u0o����U����冱��5�r������m`�o�\a<���Bۂ����}J�JT�1�~J� X�R=�oa�|�ꖹ�W���������8��v��u�]��j����Eu ��Sjv�Q:��`\��8i��[3�*Y�W8���tי��� ��n$
syW³d/~h�,�m�H�aG�����g�a��Äd	��ܕc�Zv��|�ѯ���S({NO���?�+�%���oʝ�\�[V}��\-3m͏����w�ȃ39�d�~p=��(=���y��Xt�YN3.��9d@r�u^S	<��e�8�'�i��KZ~�t�|�8Q6.�F�37ҡt��a;3v�Ό���f]w:��%	l�ݦ��{`+!+�/�o�{��o�=K��J��@��tP�� E�p����x�=�.���<kX̕$�kd�B8�Yª��ȗ��pn��~D��i��|��M�����y����9����[�x#���apޡzk�p�B�q�䓘ʒxq�摙�II��y\��C-H"��~�I���]�P�QUK6���kh�������풛	v��&>T��|��tN�����)P/}�Sz���UB�h����(X��F!�C��?�ǔ�4����&��SI9{d�k���F�=2�g6.�fL���k���=��n�ۺf�� ����ʌ�+S7f,B�YB����m���f3(���F@ypch��� �?T?�۔8zm��Q"�����|����;,��,z��³���I�}�����%?�����!�x�2�c=��&=��fr7�E�3�P!p�]e���$	iX(�W{�x�$�M�^]2�oY`n(�X���l
�8|�Z�:�)n���e���2"1Wj$�ړ�ҜK䇅mh��!���"����r�lޡLh�)�շ�>s���8S��7���W"�3+L�<��;�����5��1�(9���riR�l3BW�e	���4*zęx�V����7�,�X���y?�*��>��^�;=}��M�,j\����갢�c�G���c����c�;~nl8��Rf���_��q�ة?��f7pә�0r�A�x�]���?��,}�ѪC�����$��;��:�/!��7��rk��y3�8E��%[z��b�1`1�}�9_LKb7��{Sݪ2p\�4�<0�ٮXF$�|>�����/��S����a�0����S�g�;=����p��\\j�+e�+_c��F�,ܪ�4�6<<�I ==��|��ٯ��W�o���Y�ԃu��S��w�����C��/%�l�3/�]�ѝ� �~Y@�#B6'�ȹb��PC<���s,�Q�q��w�(g��Z)��/#�~��+r���$	�+�Y�9OT�h�h���]m32�~#M&����"�U�HU!�g�uft��SD.��/OpIHH�Z �v*ߒ�U6�~�W;x,?bOU �&����(���H���!�qx�P��bš,n�(�h���c���
�(Q����\h�����G!��3pH�o)�X}V�>{l?���z��dB7c ��A��AG���/ j�:̩ng��-tf�p��Bx?K��K�Z ���
�ރ����q�1�`�cd���?�.y�ϴÙe������ ���6U�s���b�tx�ҥ�..� ��7�xO��=4]^��ObX����2q��mp����J����o�)/=-����f�~�?ȃ�/d\��h� �ӱ�Ojv��&�ȑ?�UCW�Źn�i<T0X�������w��X��sag�t,�ΐ��t�����u�uXj�5t�N)�XB�mB�
�eY�IU
��tz��v}�������GC\��ĭ���\*y�����?�����9~T�g��̖H7.���4A�`�b#7�4"
�`��p^�Ҽ�p������x����kgK�Gvv
��٣��+�ڛkK�!3�{^���&{^\�^Ž�������~�����<�3��u�Ё �.Ej���y&r)s��_�w�Ȼ_�I}���g�� |@p�m���}�ƞ!�9�=�ܚgu�M���w��i�/���b��F�܃8-���?���5-A�̷��w=Rz?տ��c�!��IoVP<��ޟ����Ūb���{q�"X�R����6�f=]�f���uTi��yCq�POZ�1����/���	�q�۬2�K[k��W~|�(y�I��������p�>E$u��vJ!D�o�猅	_��?vEw����[sgb�2
��֝��̭%��݂�4�\�Gy�AIOXM(E=$j�-�$�w�4�����Kj���;�^�P�۱�R�����e�Ֆ!g$�~���^�`�K�[��
��S�|��'e�3߲���T�:r�>Rm��iyG=�.]x�R0$���e�������ڂ����X�Nֿ+�JIN.l��aD�E���g���N��֣�ݖ�ɂ�G�o�+����]>��AF�2� 1�ެ��oF��������]�Ѕ�)���8���5'CM�x����\���Af�v�tY�s��[��F�ɪ�B��O�.$g����C$Hp�ő��R������(�6Q�9�Y)�����-uk��jg�l�ܿ�P��Vyg��3x����y`�Iv.��=���AJ�Cj�j/r��JĦ��c\�ε�bjdԸ��m�wcǺBLZN����]�,��[�?�<��~��J�V:�sR���{e�? �G������p���!���j�����V2�߰C91(����;1�̂���y6
,w=锔|(��!=Z��{e��@�O��6���AӇC�l�ec��ם8�
 P�s"$��I��F-��#��2��~j<�q__�V�{�:]Q�Ś?�����i�y���7���?��6ȕ�|_v-T7U}ٕ���������eO��,���<?��e��G?����%��G4a|ҘHԓ��>$�x��vaۍ���4k	��/;�m�����؏��^��)������j��=ٵ`�59�����"^���i��$o?�[���X[s�5;�Z�f.��/Pe�La�\��x0�\c���8\�15oM XR"�U!�/����0�+m�Z?�~����udtƥ�у��Q�\&�!��i�{���t;Jˑ���Ia�tҝ碘�>M6n�g1����L�&���l�m�b2Go�WH���֦��/@�z��O�&N�)��J�dHj����Z���hs�:����v[��t�uN�i��W�� Q�4����;�>��z��w:_��:���?�2��*Q
�er�c�*��;�~\���%���ҝ�
��2���:D�dk$��6������[zX�"���GּD����pt�5/7����5b1�~=��C�C}e.]��6��sɘۛc]QZ��k��=�(����MHM�i.OT-�^����>�O�QE��=�@�wd���H�^!�&=*�]�
�\�ꡒ� ��\�YB*�	�];�H�m6S�:��܌Z�SLt�/0n�n�g4_��Vs`?�w+����	۰��%���J/�~�s��` �{9ó�,ϴ��FJu����d�w�|TG����7>8��f�]��%��tD0
�lJ�q�����g0����!/nnO�mj�N���L?�t�ŀZ���utuVwa���k�w��=�5안����xl^Vd�<	�"���e�󖖵�,��Qv7�m1�щ��-b8�5
5��O�OB�Bv5�ɾ�务��Zd��	ɟ���!2��������))ZW�T���1���Mؽfb���G�'Yr��v9��ݭ���/?��;3FѸpg�j��5"4Bv1fC��c��)�?��\�!����y���6,�u+��y��� ,�f��Rǽ(��N��UD.�I�:��)_��a���(�;2}�6�A,eٳ&s��Vh����`�A�|���(I��j�~y��E�\�[<��k3]?�E�<Œ�B^�����k�T�tp��	3����+H���ױ˫�v�*@�E�/-`2E�5����h�ǈ5�і$����Xk���}�V>P���D`ȋ�"Y��[���/��	^�:QhRA�l/�B��Ƣ+��~A;	��T�yt�"��g6E��9����*Sx�+/N�)i��@�� �9�Z���� ߐc��%�eW�m����,����ڗ�b�!)��QI���#�ѷrccDF�����G
4+B!�&�*I����*��k�~���-�'���rVƝ�O�]��\�8��)%���������]�U�� �tv6�U��)H���o�#6� 7��Ⱂe0�X�2�s�zR���Hf�]��+\W~l��N���?ՒS�	�|w�����`�]۵Ӏ�Vh~��@#d�#�ʘ[آK�����t�Re�'/(�hƭe����<5�>1�y��%n��s��ڽe�|?���&R|T����S�B���#]��C����$�~Cܱ�B�2�	�7������nv����&QT�=?���{��I���s�0�Ȣ�2y���|�w+ �*��#�'�K;��wٶ�A:�AZ���Zr���AJ�q��A��_�z4%�Ys���VR�ְ{�T����9��K޷ɜD4kN��Mb�$ݶ�<�B�W�G�g[�VUQ�ܓ����J�d&G�WǸx�a�6Al��=�d=*{���G0��F��ܰd����������}�U� ^*���XBj璁����'�/���n��^��M����t2j��J��G���j��_Fm�ej�)
��@�>&Ў~�#m�u�WgR�{s~���G�	��b��켿7 ���?}D����7b�N��vI=���Ҟ*j%cR�-�6
��d�P{a��Ǵu����1H��cE2�m���_S�zU��Tu�زa������
�j���А�	����T��ct���k|J�����#�R;��ޣ�B@7
���lz�A��K�\L~.��^kx8-V
��n���0�F����0��%1�,
7&��i-C^P2W2C��:HV����1�)9P�-���Ù�}T�LVC�[V�Z�X�}�a��/̇&�U%qߋ������ݠH���6���)8t���թ>* ���u3j���e�m�!Y���%�;m�A^�.aS�Dig����_e�#�ƅ��@������_:L7d��~��D��O���s�iä���a��"���X߬�=J���Y̤٥?���I��!W��|�
 ��C�u�/e���4.���R2�~D�S���0��e�m�>�zd�uX����,4��k��<ّ�����=���L��T>P��L'0��P	�RZMԩ��q�%��%> ͪl:X;��*&����!�D�sA|{�k�9�J�d�7���7�����-E��m�Io0�����"����G ݜ����
�S_�W�� K��k��E���.1��_Ǹ��<�u����O�QQ�O��,�U=>�E_>��n��W!�v�OgF�2�����b�����А:+�v(���#[[���
uq�j�:&��e����#���j$#q#k�lG�1��Y���]�N�2!;;{w��U��~��]a�G����A�DN���4thl�J(�o�������\��,B��a}�<���ч�DXT�>J��C&�K${>���g�V���&�$�K�o;f9�N+��0��r����T��Xfy��h�X� w/�I��_�'���/��K222S"���cL)=�<�l��7���o]^�'K
͊�g��Q`j�����X{h��p#��G�i��5����H����C�ב�;�h��v�C۵ٙ��I�C���Y���>��-�r���)#�����-���F=�����r}��
e]Z������C����BN�S


:�$����	a�{������'Fa�Mu�G���7p����Q.���D2����#�#TxM-g�״?�&=~���%�A�k�i�ܲ�h���Q��VB��l�O2N^��E^+��>��D(���i�OXJ���`���@����~O�n[�G�a��K_��"w�������WO���;]�� �+�v����;�T�A�+�9�^=:k$R���UOl?��IP�� ��w��Ժj�D�;i��>�˰�LKQ�`�0O�i¢�`�� ��R�M�gɞ�M��m��W�/jʲD�o��Ny&��H<8%Zl��6�|a���,��������j@�0����<?��KD�C��w��/�GM���T��t��?os�=�"_��ĳ����S�!�����D��(ԥ4�K���o7�� �k�"�Y�Y�Ģz�pN�[�ޝ�Y
P>ftG����}�ݨ�l4�{E��:> e��T����dT&��c>�U��`��{ޏN��
��T5<� \27MM�☀Mϣ'�����������B�z�S���l�A|Ǒ�`�z~�
Q���
l�ހ�[�+7��'��l���B���DN������4�0ݽآ_.p{���+�;�ϛ�끕��1�'��d��eg�뙚hI��cG]N���ͯ)G�A�����p��:��كҋ���P"N��/6�L�C5���s�oIO�X�.~��+�j��� D�ġ$-2��Z�Ws5��Ni,-�>���lIҭ#��w<������rz#�$6% �M.C�xSs�r�ݩ�AZB�%f�N��4�.P��8�A���!/����sx���-�[�4��XV<W�u�`���n�KΌ\�!PX6���՗�.���.F�	�\�\�[u���|��`�4�^k"��Co�,����د�,}���|o����.2H�j,quoϹyh��?@�'r*�6�����-���P�7<���/����ˈ�o�~"q��EB��;��(V�;]���z�S�M���w;\�F�*������B}fu^p�# Q߿}�,��Sqe��n���@�̞<~H���~H�c;%d�R������`��\Rўd�h��j��|��N�UVg���@a������c�3���!�c`kck�ʺv�����2dN��hW���"�F6���<�'��\����������Bb&��������G�-(��[���RXʐ�#�����0Dsٹ���& H=q �ek�;'j?}�ob�u�5��:��A���q�#>�� .�����@��IY�� �Hz�f�m���I�E�%��Į������� Q�+��9���%S� ��A��:%��!n�F6f�� �ϡ����K��T��5����8���_!M�#�>�;�����eT��%�G��fX0�J�?CNJ>5&��HL��@%=NG�7�=H������yH�>��I4�ݽ�`�YJ{
��l��>��2���N}7� <���h��![��Ģ`���S`��t|<V�F�ܕ������V���a��x�90�%M�Z�7���v���=;��x!L?`��>�y��i�?��C���P������2Q�{���[�.��dN�q�I2��{�C�_nw�Di3���_����hj|]4��3z�V�a���i�\�Z��߸%������}��=�9ee�}�'sK�1���sP��|>�^j.!˵�7o,�����/���6��A�v����O{�� �U"���U_>��~��@�n����>����-E��ep��!_K����r��M]�ʁ~��T�{U}Q�3M�^��;	w�t'�߀�y�y�|7��F������C�x9��������>���vl[5-�N>�*�+���p"w��9)l������6�{mY�Vq��Qߙ$HqB���o�^��+���]��Kl��ݐ@�����Z<�Z7�X}{!��]G��fxY&TR�J�K>�G9���+Z�b\ۻhIC��� �,�R�)�S�����@�9�D ��R�a�!J]&�4�l�w*H=5pg���S3��h��D̗<T� ��ΞS��%�4�����
�$} �H�����d����)�l(O�Ċ,C\av�7�GϏ�v,��g��cP��>���"�!�M�7Ӻ��r@!�̳[/R=BB
��JO��{=l�>�C�ͩ��eC9�M�ϬF�ZicB��pT�ˡ����%�����o�%����[MM����a�A���l��F
hm��֠�h*r�4Q�I���F8�3TFF�1�|���W�P��鮕G��͊�L˝�D�V-��J�HIn��Ǵq-�J�����h�i��,����k��S0���@
��݃ƪ� �P��Y��U��1���ӼG$�1���,:��V�\>���BWr�g�F -�{K�M{_Q��.�:%��utP��p��G��9XG6DxEة-��Tk��xIrY�&�d�Qnڧ�|�٧n���|���N%�/ޠ�e=_�RnR������Y�����#q�͆�Y�_��_��Jt=���Hy�=�b�r��yv{-���w�i��[0)�7K���5B1�1���7ba��9�۲L�%��F5�AJA;�2<��^%%%<���w� ���'agi��9ڰ�e_~�?<���APT&�k��Ml:N�#_�+�脭3ğ�-��Z�cv>�?z�ȶ�ް�?p��fJ-���������T�\*N��Tݷz�U�m��J=r��]�-�Bg~��'H�,qR�Cg(���_=��������5������u�)�v��5o�4db���m�������ùx���J~\�U��!�-C�����+���'��䠩׫6�RV��T0��S�31�d� >����S�!����;;U_�E���C�>`��f�z�t/+٥W��&񵓹���-��%41#4�{Myi�`ڙ��ECS�漸p��;���IN����B�"��q��+e�a�����@��� �!g9��qQ�+Ԃ��<��pz>�L�z˕��7o�#���v{W�4����U�Y����\��#UD��g弟'a�U���9XrR<;��6~W�7�Mx��p�E��<�>-dTܺ8Nh�Ĳ��h�&�E���+sT�.`�g���K!�͢;p�(Dg��W���L:b/ĖG� `�W���#)�.-nk6=���Zj1�4��EN{E�s0·1�P�E��]�oSd��z@4Q(�Z"�ص���'Z}ĺMѓ�k��ſ��b�$qL�u+m��[*b�6��T�}�s\'�uF,��D�N$����Is��[��H�qS��i"	�h��m�G2R�oK#b��|�%��k{���x����yNz$mS.��3����ݮ��X����M��!I��I�F���K��lA,��X��K�4�w-传��Ԟ�C����2�}�Y��=b��Z|Z�J�[��@���LU�2�hyl_Uh.1y�Υ�:K@
r�8e~a!�
E��ǒ��P�` @�Tte.=�V�-7a}ҿ�\��ǒ�'�o\30��r��Hn|���C���I%�k��jN�V�G�����Uﳇ¬�{}��`��m������>�����A{�8=8;�!�z��݄��r�x'<m��&l���VI��U#p/�9X�▘� ߨe��}!`������b�l�8hL����1�f��(6rt�S͌f�+�i��^k��i_�b�7��]6�@��@ͧ��ӧ��l����;�������	�KI��iY۶����:���]?�.�v���oiyRG��S��NPw>��F3�B��#`>���
��b�4�@ �f��n^AT"1������3�n$j�4�#�~������N|�?�E�7-E�5�fG��4���=$����ܾ�6�54�'�˖kiݥM������l��ƅ���T���y�!^��7zc.�!�.�Z�-���.ʔJ�ST��jʅ3tl���R؎`��"������G ��=�ݲs�Q>�UA�U�Z̶�^��m�^<o�{�H��೉���l�����폎i��h�.49�O3r*0��m�v�k����\#2�W2و��b��/T)��v��Z�?s��v�X�X�1���G�÷biZY����}į���X,� -���q��jr�j<��ߩ9��ޝ[z��T�ݽ7��E��`�HM�
=A�b��rp�q�ω���>�Z茻*#h��p�XU'h��y;�2�t9��������Y���;��V��E0)s�[�����B��Ǿ/i�BOZ��3�%yAp��Ϊ+��p�;�׻��'H
��Hp�eg����G�g��$J�u�+��k�^K�˧]�l��~� qE�̢��5����װ~�ϟ��¸�C�%�FH�6�r'h�z��{m�JJwW�Tك��{n�O������i��46S b	-�;V{��!�nK"1ʱ8pL^�5�\�B��	�#|�h>�;�8 -/���9^+A_'IZ�߀SI'��ML�-׍���bZ�z�^Hp� �9�ɲd����Aߥ��~�Y(��6�T��N��`�^���#E��R!�Mn'7k�=(?�P1_{v39���o�&�,*[🗔��%�m��MCČ�F<������:�F,�*���"1�J!�=��l{b���0��09@���y�9�Ka�A���.�d��/T�f��� ��R�j�
M9>�ҝ��:w�ו_��`|"1ߵ�6w���8��sn��R��pӅ���4�۝���	�\>xg���f[x�L6�p��|ͧ4��A5�i��]ʹ�y4w�Im�y(��>�by��K���Z4 v`��(i��܏�ʆ*~P,IF_����wfe��S��jp����j����a��`���:��Ҿ����nd��M_��]M5�F���<p¡K�Y�M��Lyej�}�p8x�[���yl�{j%��l*��냤55���C��}7C�k~��\XѼ�6�6r��翞�h]g�se�n5d�� `<i�{��(���2,7��6������J"�Ώ FcKޙ�H��� Q�͒�T	0�Րa�~�wu�[JI��3�W=|F� k�I:TC��Am����γ ��f�끞�����><T�#��L���I=o����_�8#ڴ��ـ+GaU�x��2o��ґ��SqNn%��6Eu�\�G5�_-}�_Y��L������e��v����� �6� ` ̔b�;�+�A����U@\:z�@Gװ��q��r8^7��#y_zX�i$�W9�-�������T��K飒��m˕1��Hhu`$P�&[}ҪX����Y]�p��u��VoѼ���I`�-�ݮ��`	�����w�*��X~� b�n���K��f��RCHeg�%o p>E7����m�����$��V��bv��ݢ����]��}C���0��V+h�OYn2m� �_�1-W��&-�a<*;�2~����H�����ۑ0��\�5ǖ��y�ھ��.�嬶w+-�ۅ���r����L����*-DN)G�#��oВ�A#�����u��^�L����FB�ru]t��ww�nߎ��o��8�����6ޖ���!�nM�[�s#���*�D-<KML�s�P�4���~�;[�
�t��$����F؇=��؞���kԣ���o�҆��z�~O��C켟�]��o�$z&�Ǩ�}+"�Z����7,�,��4�ߗ��|k�V������>���΁��\ᾎْ�]��Mƙ#Щ��_۴w,v�"�(����l��Ӱ<�F&�����y/��/~�[�_� 󗴥/
��M�?=��Q��kt�5F̩����NE<��]�@����,#|��ȱ�fm^�K�U��%J���(V�?��y�ȩzmՎfG&��r��R}��ITt~�$"�bz$�$}��'+*<��e�i� l�{��L6xq(v�Y3�ش��;�|KC�e�㛪{ľ�\e\�_�ݣ�T/�@��[��3��>�/~��VA�����93k7Z�h��l�kx2}�ưkG�ĽGjg�9��`Y��uG�L��!FZ���֚��ޭy���z�e��f��Y\1(=��)ȃ��#a.V�r��>�$g�(��ة�� tzn�d���;?OgW>]J���jD���3���#~A�wD�u����W���E{S��e���[�y�N{��/��Z�q2�=2�� ǔ�:ܽR�Ihdb�ii�0�xE���	��mִ�.⸥0{���f���;([�)����������1��[*��1v.	�6�H��)�hg���9��}�N���^�`�������9�č?�ZːͽL�T��X��ϳ�}F�-
�ONo����r�dj�֙�LWgmJH^�	��|�m�����Q�������e7IZ�k�]և9HGiH��}=�b��-5��_��YP�	yC	�D��0�-���rI�ݲ u(*����S(J���͍����W�nf7��71��ٝ�)7s��ןp�gBhNNWծ��RБXK��}
U�C2�����VI��Ƚ_��|1�����Nv�*ŗT�a�:�'�
I��p��灕�<�"Ku�OL�E����� �-Ub��Сz���X$6�ml�EF���ޒ��j�2��������[O�flom���Zm;~5̛�d������?��6`��l�M�Y���%8��s\�:%Z���<#\�߇ޒ,���ڎuuZ��ߍ@wr�9����s^y?_��i��#��G��8NR��?J�L�v�,�b�Re�*_��a�M���5نr�����%W�B
hB���"5�D��C|n*��l:���BYSY8>�_T��i't�8����)0������>��e��A-���f0A���5g�z���h	Ks>$z�ey���f��+�ɮ����}"�d��B@b�9#cgA�39�{���Kͼ��L�s.a�9�Q!��������@GF�΂��2hn����<]�0w�'����&�-�	o���l��**�<��ⲡ����ZɁ��5l���t��H����/R�Kj�9.�/���Y�����2�p��>��
�8k���*'.n�~~�RU9�K��KO{0�6P
.p�R�Y��{�5[�l9Tc�8|H����}��G�_YRWy�ߙ�B �R��*B��|��Z?���vn��KU�r��2�Mvh�P��Ѷ�T��"I�߾[���x^����zȇ�ծ�5	��u�G���*�нy�n؋�H\���E�5��H "=���l�7� ����B��+I�f��8�.�$^��Qy��b.zW�O�};��d��'�P��܆E�i�E_?�� �+X˿��(>w>Z�E9�P�V�����(
��r������ ���0�!u8s-9��N��+]	Lg:{F�RT��va�s��&!0�_j��O�&�DDiZ��5u��u��=K�<̏��n��� +�ܼ�ڑU�?]��*Ds^5��:�r�j,�ibŵE��'m�.vn�~7u� �i?wL2��Er�/M������(�k�P�9�Gj���|rT�ms����`p�S�%�լ��?d��^|��d��fds��u��(�Цw��k����x�Nw��d��=u�2P&�
u�󡙴���W;�ş��J�}�&���Ѝ�c�V�z�-��\]��:���؈LT���}`o�"�����Q�+Q�ҫ�	ټ����q���N P�R���n�����(2$?^��ۛ���#� ��xs3^be�Ƒ�Lg}�Q�(���S�X�n9�\�vԨ\*T�j`���r�"/�~8�f�N�f"����LN��������=�d�����b��`*��d
"n��BaC����Ԗ�H�w&��t���<i��Z�Z
�(V�"�*�ퟘ�sBSRR�����6�%AG�s��%v��cv6����@o��^f���>��B�
��z0���\�� xtW06����n�]�u����pwpy�5?pJjB͖~<��d�i�4��?��1�{=cC�����wX u&W�ұ�q%|2��_�q��8�-EaZ~�O[���E��Ēs�x����v��ز���E�g�����X%+�euY2!ĂCW�~+Hl3���̯|ev���A8���ٯ�.�}=	�* [jH͆��2w�PrH�=��o٤�����ƱWCuC�������&~�+jٸ���H�TI�'�d-ͿTK)_W��)�WE}�:�Gb5G���W%H{�jK���0���k�{Q���+���	3y�cz�y���D8zV��Rn��Pn�ҧ\���K�j�+�R����&*&W�B^�ɒ�Qr�)䥁߂���W��_�Ħ��;���'�|OEE��{��nwJ�~�),�n�V/R��%���;���o�.��?{�p*���.��/��B?�u�̎�D\�_}�J�dU�����N��+��B��'@Q3)��5u�c��\�r��6o{hI3�PN�e2��>8�촳�s���
�/Y«�*|]]l�9t�Pܨ�'3�Њi7�F#���^�į�KKf��'�h@�$��yG6���VNP��}-Ԁ�n��\X�^����s�ph!"�2~�۝�d`�Fݎ�<kw�w���1# �p��M�O}1�GF�A�Q��VuϿ�/��+�)f�t/�����kӺ�������~_bWv�v�:�����^O�~�_m�_Ҳ"��!{�� f��-��mB	���5��|q����~��x��}%�Y?a��33����Y=ys��9�ސ4O�t�S�G%A_���U��� �@ʘ�ћZ�������������0�� 2����� ~1|Vh:��T�*M�Q�S�7��M����k���K̈KW�䪒.Kr���t���O����6����Yw����><�#V�	�J���<{ndj#�.א���q��jK`���Qt���n�7�T���3�[�E�
�X#�~�z[� �()M�@U-�����[�XUD�ER̂�!]r���w�l�Cݯ6o���
^�����ǈF70�"����P ��?{H����fn��N�d,���{0��ji�N�������$��BikW��|���C��4��]��.�����5C��{Y��)�0-*�M'џ�Itm���J8�݇�v����i�PRy���KW���B�V�u-�8:�`mf�f��_=6GI(J�bv�8��z?��׋[������C��Eo�IZ�����pͯb�e��Vf�_���HJ3������Uj�0��6~X�z
o��]Е7Q7R{Ɲ\��G@�D����]�{�^@f�/�o�k#�r9��cI|����E��oȯ�6�Lq����kҤ����\m�E�R9�@�j�͸$+Ѓ|cΊ�)�L{S���|��V%͚k����{+��Pw\6��6z/j�i���,vѼׇb�;�Gn�s%�c]�S���7�趖 �GD�	jNF���F�dO�N�g|wVN�~��|��H�
Ġ ���!N��l٨����� �s5U,�d+R��Q������A�X���2�f���o���l���`����hM����'p�e=z���\��k��k^�k�CA�A��+�^�{>���M����f�0%�uWK�ȿ�(�UR"x��N����DJM�
r0:SaU���:��a^�(�W`��_����/����A[�N	o��-|���~��P��moq�I:���4�|�/���w�J�s�z��tW/q�H~���_��2�`T��m`�fs�;�*&�tMÑ���Ĕ�I���
����_¯��A!���w�m�:�����ڿ�.Re�t����wD?Ɗ�.��ӳ��9� {���13��G�٘	������5��x�F�����T�"�M�,�i�O�o��y�9�����J;k��7~fT�5JGa�Ե��uB�߭�T��w��/�+�'Q>v������e?t!��U��Ok.۫��Ҩ��5J ՙ��>�<cp槜�"��z�n�)�1P�\��Ҁ����m�Gt��E��|M�{��*8����V�Bz܉�/pxH�d:��� M*��uD���8�̓��� N�ƆR�"N�L����;z�-i��ŔEI�{�N��l.H;�D<�\�}k/�hi�a�ۜ5_1���yw�N��h;Ţ�zܜ�
�xQ<�}l>x��^tK�[J9������a�lT�+�����.���'_��.�F��/s��Ϛ_�y��c��X��f��FD���)	�ŭH>�T/`o�y9ڗ!lfh�g�~@顯c��U�m�䫽�������*y�;&!	/�m��-l�rľ��:���_q���H_�r��Q�%k�Eާ	݇��D��������pQ2�;Ý�&��I0V[u���}(�L��޶�
�N�ɬژ�O%?˓�
mӒ�܌� +L�wg���|$z2�g�ø�$��J��.��&���p"�(^�^Ψ�Lf�Z�9\�����M�B�F& �\�=�"�X;�)��:�f��2�YB���ފ�4�m��V�D2S��.��7,!o�;}��������l
!�
s�:�?6�٭�/�;�5u��J�%��#�?��e�]�uH�$ecs�5ÅmFk��"-�����_x$B:���Z��6�.D0WE�Y�,M�M�H��4�+���g��c��NDMja�����8��(���ှX�����^(X8E5��D��v�*�?��{������t�s�~cqzg7��Gc�@���!���ʈ�N�@6K�	%f���{ۢ�i=�A/iZ��SA���0���>����K\X1rأd�[��0$��S=w+c�����䏥<�Op���_F�p}M-cf�˕���ϻS��r���F��Ү�z���;o�,+��.@�*��(QRP�=�3Y��`�\�hy�H����>��ԲZ�S?;W�D���MTk����rC����������Y�	�����8h!��mG+_"�,R��<T@�������鵹?A0J��|E���B�%��h)Ym/&��z�~�¼?d�Fz`g��%F�#�wg�E%�[$�(7׹
5�)�t�ɜ�O)�6}��T��e��*��E��ܽ�]N�Ubx�P�[j�y�g{��J�0+2�r���c;ع(�#�r#N�u[&ȡ�UzC)~d�	~��SL���\�_Ͳ�9���N7���i����T2�]w�bj[G/�/�'���E�������� 6�0���߽u�X����1�����H�Tʄ�vf�v�=���u��Jo
��~9n"�l��^^W���StoG���R�KU9K�PN��ʣM�+�FY_���yȞpi֝J�a �llX����
ꬅ!��R�ր���[�}ZTm���jؑU2$ǻ��[1@�=�K��� �n����Z��ї��)@w�����;��7��lȵ9)�V�,���h��Z�7����ߛ���	��������?�l;g�Z����3D���so{�2�1�ƈ^��o��+<���KOO���HsxdB�v�mrhЃ.�ͯ��lE;�9�J|�u�V
;��?�\��G������)B\,'�T	�{b���U��PR��_�u��X���:%e@7܃q�W��{+Py�R���O.z(a#q�o��l��a5raX�UxP륖xP"�)s���:��m�E0��gA�jg_��[I����o��iԔD��H/�DP���^�pK������|�d
˚�&���@��N+2Ōi�v��>gj��c�v�N|H�X���J�p��\��?�����!��d�4����}k1a�����r��X����ͦN���6(�n�Q����}�)�i����g���熐���ʌfu��wΖ�wȚg|;��}jbz���ڜ�.�O����Y1��7��c_A�,0Uͮ�f�h�E`\<��z<zo��qa�'����]��W{C�\|�K>�o��t��C@FO�l���^wAs�!U0?��:�*x�1����c�ڽ����!c��>K1�Ξ1=���oul���!D����� �fԣ9Pj٥{����8�0O�6�J���� 7[Q�C�v�&�������;)��T�j�<�"����V�6����w9�>��>WT��y��),�=��
J���
�%'_��Yw�).��y�q�6N�OS�8���!��rt3�/�\j�GKV����-vg.́�K��p�FC��e�&�'�<�t6K�G�v�0�[�9��������"�6�W������4-�T �J�G��Ά�6��>��e���/���vdٙh�)а�v��d��y�L�U��z4�q�_S:sK��\��É<��\��WWjc�����0=t]��x��e�VEi���0�q�c������y���F�����Ұʏ=M���Ģs���|c*�)o�rL�(����'�X㸿��?��g �D�CTm�J�4(�0 � H72��� -]ҍCKHݢ��1tw8t�C�}�s�_���j�{�[��t.�0���u�hc��\���CW�EJ��!!'��t��Cf�Zk���S���z���aZ�b����c�4��qA����8���/�G2�I]f"^�	�q�}EL�� E�f����W����T�Ӽi�	=�������,�S��/���=�'7�O���Q��*4W؉���ӊ�ʻ/�ء}S�o�n�\5]�*��f�-�F?�5
y��#^=���������	ŋ[��5SP)�F��1���7���<���T��ؤ�|jm����󂨁���f,��Z�_���>�l(�i��'Q9�p�i�嫠y�Vc({D�+�OA~nhQ��|qhR�^�P��˲eiTߚ����3Ґ����� /B��C{Re�:��vGUBޠ�}Ǿ���z��7a��>�(��WL��E���*$-
������=i7��u��[�]���^��ڣFU�1�u���kdς["g1��ϗ�;e�ή	�贒Q���p%�u�̥aP1}%a�6Cl1ðSr8�*�%��	�Ǥ��N.�M$�߿����l�.~�j|s|�U�m�<�s�o�^Kф<�;�'�LX)v���/�tٮK�F0Vx+���v�]s�dk��,��bm�i���R��������TS��P$i��{4�Y�X�}Tj0��m��|��Im^`sxS��]8Yg�鎯��>k�o�=~���8��k'i�ʷ�]��L��~��ޯ|L���a�+�"ȱ�:�ފ~��X���X��Rˏ"}�Z�h�0}{�v�I�ȃ��R�=Ks'R�����)LK{5��?�~J���?� JX�٧�G�����ړ&�<N4�,���,���9k��|�Oc�߬g�x������,���<ਅ�Ϧv�qF�!���������	&/��3���:&u���}|�\���3���R>���N�"�wV7^�Q��"K?�Z	~w^�;�{
Bd�$������s=<4�"'����@���P�n�&*�B�k��y�;JV�b�c��������
��ҌE����Py�A�W����w���+�}	p����	^_OX>+9j�w̻�܈�v�eH��t�q;�磅�S�O��M��
�qys�ss}��d3�o�]j�л3U� �Nї��xo��(U���g��}j)7n'�=>G���+**6��:��h%���{���I2�۔ٜ��-Vi[��<��p0�u�K-�X�Y��
�"�!F�O�叇Ȝ���uX�Zt��T!D�.t�4���-�p>��U�F<49Ibb��]T����*�9�_����?� ���[�F�y�ġ������(��N��s������ݜ0,uO,p�?��&qh��k�K|e�G�#r8���oL���Z�k��9���4��2��d�����Ԯ숚hmR����������(���o8���Դ��4�bj����~X�쇷��^��)�}m�����Ϫs�4;��:�2�.��*��3��}..�A�=0�}�}���]�?	ԏ�e�+����>F��	���y�BZ�kvh\@N?+Z���Sn)�V�-��ä�\t�Γ�M��|Hy�}+s�5�g=/=)G�`�<�s㷌��`,����3�g�!����n���>6v��]~��;:�c~p�'�ebv�>�(M�c�2�b���~�A.s�5��z#r�l�`a}�ZK�|�Z��G5w-#��K���Q�����>��>/��j{����O����&����e����Eh�Q;�I\*��שR�qq�,�6j���0���6�!W�p[�����P�.�2E$�Vr?ٗ�åv�fL;�>;���R����Ȝ�ƆJ5���Ƞܛ�؃�p��ʛ�4�X*����@��::����C����k�؞ާ���]��*AG� g�<"�F�_{��r�|���HJ+��a�߭�=*^�����C�t�ܯ���9��_�d��V�[�Dt��!P���b�+��}��ϼW�I����ZsYg=g�]+�Kh�N�S���n��}��$��b��_Ln�2���9�Py��T�L�-���\�gu��N�ο����rr��ި.�G�9����o��{�r`@��4:e)I*3�����+EѸ�dw}ï��p�-��l�w�6��&:�r7F���4�ִb�g�:GrJ^��)�5�1��
��2yVD����=���e7)a]F�`SD9`��L�Js�dW��N�����9Ɏ*p}�a�����!8ي��������*��{�k�K�B7���`�諍����)�ic� �݃gm����z<[snq�54����/I�_��ˑ?�>N�}8:���]���uK������َ�u;a\�2N��Gdx���O���ʂ��>┚�+���D�G��ז��� ���|'�����g"��Dzc�g]�e��L�nK׹od�*��T�|<�kҩk+า i|�f��8�i�-H��=��2����E�U�#�*�FH֨�ɣ4��b���}�ӏ�������|�U]�fSC�c�+v���c9�@��>T_�1v�:<���,D���ƔG��z�ʆ���=aP��Y�l�le�
o$���>�N�N?�N~p��*O|�@�@��_�����=124��Z@}�p��R���_C�g��M���OJ���E�5�>�O���Ƙ3)���VvM����<���7��DE�v}ڵ�i�$m�C��RG�4�R�����*�u���/���PY�:��"_�Y������?���-�[!:^�f�����ArH@ ��l@�g�X��U$
viA�/Lm+L�S>u$�W3ֿ&�Y�otf� ];�]�����_Qnx~����;�ո����I�ܜ�Z�p���w�y��wp��|�pI%E0��\o+?)_�gZ��w$�0Ɂ*��z�������z��N�'� ��8���~�/���Pd��G�i�d��$6�]Yul�����f�j��v}nӴ*�, fuKP�i���4�W�w�����2v��[��A�B���w��2�".x�B�Lݹ�>�jiC��ࡸw��~�ˢY��̝.��C�eY�����ZS,������'*�Ƀ�`�;�Ư�IB
��8��34��w�M�>Ф����ٵ;�\�u������+��C�Q �|�oe��Ðy&��#_�����4��R��ݑ^+sW,�$��W�K��&��/x\L��찂\�̍-քX$�����L��F�ꐊQ3DW����/��{>2� ?���_q�N�G��U�NA�$��a��}e�ri�o�3���g�I<��&\��ëY�?Guj�(�4�����w&���z;7U�DlT��a���Be���mk)��׋;R�N./	�t������X��hNg?�a7�9M�g-RTf�?�����V��l�>��ĵ�Tҗ�)�6EǛ�6�'!(�)RyϠ�̚��?�� �	1�s$��ir�
~|t	�e4���
��c�	�&�l&�D���*	BV��4�x>.�]�8��p��4�!YW�l��3�L���E��,��;�Kb]�g��,�#���ـ��h#=Z��rSԦk�輁�n��['[Bƭ����sDf�ܫ�G(���7��W.��sf��&��e��~�*#n���uD&g�'����!U�4ý}w9���ڨ�v��b�쥫�m����`��a��:m��l�Iѝ��lR��Zī��,߼e3�w1��jmK���$c�!�sV�7�_FIcʘ��l�~�$��	E<�`C}�;�Έ������.�R�/���"��r� ���m�oJ�Zl$�+���[f�x�>QJ��?��<l/.�<����:� 3S7:�>�`�(�5�d�Tx�a���UZ��w"�����x��(3e����ەdbT/Qԇ������v��i~��&˹�~��m�Hϸ������D����J��T������2���T9r��[ʪV����8Ȳ���v��&������Z��2hO���Zm�*,,}��{%s���������.`�,���y��@�ʮ+l�~�5�x��Ĩ��E�fE�2�D���g��[���9R�gN�8�j�
�D�������^�Ã�}T��΀�#���ؽ1����Ƚx����q�Oޓ��,���n�
,���Ŭ{<�}����r�+w�ێ�m�(��4Ɏ�$h��(��Q�'�t��Ö�yQ:W��~q+�P���O�����֞��L�'�+:�Ώ���f�
W����j�^����x��LFM�URqZ�i2IG�{Z��|��<f�6����[�}d	q�,g�> �C�h�$�@��RH�}�%�=V�p��9�j�&���A~타�|D)F��D_�#�Q��7��5����;Ij�s���ēu��U��T=����T����� V��b#�+Iki/'O)��/�^�s�b{7����� �͖mE�1�N������w�_�)��k��V 7��}�$�܀�q\��Wo��U 4�HZُ_ue�;W�,ԋD��_�к���jϜmO���]n�{�3�������,���n;�mÛ�#8�R_�$�v�soF6%(h����6
��7�n��lb6� ����a�
+���,�;c��;2����ˈ	hԟ��*F@��&�,���90N9�+���_�=#
/�ؒ��%G*@xh$K��٠|�4�+Ƹ����K��}�� �L�F��K��f6�VPD�v�nջ�p��e9�15���Mqv>x_c7�s��j�"��(����J����Btѳh��.z�x5vW|���;s�DT��b�3��/�2Pf��HK���g�Ҙ2I$y>L�r��~����C,���YL��r��)ݚ���+�AY�X,��2�[�g�g�C�@���l6ߎR�OB���{��QO����M��{�/f..>>�ƙ�
�2�5	�V2�J�d������<�����dZ$J����,�`y��l2�޴��\a$b�&� :k`�ި��~<����b���F��}>��/�����~�
	��'�LS���n�˗�$e��JM	��9�z�/��c2���>���
�I3���ǉ?LrԦ�1�<�z� 򆳇��&B����JMq[f�zl��	��u���q\?'�� D6�m�q���A���|��x����Ww��-A�D��3l��>�=�[�@�� �vXX�??`iA6[z��\,�p��B�YX��֣�ny	L�}�R��U�O̻���X����a���Q��tw��5�}�K��yx�:�g�*e���/�f��6��2_49��/t��R�6*�f�1/�v�}�Qԋq�?����o�"4~x5�Yg(�dF@YA�K]���?�*�������	rZ��ֳ-��;v��:}9�m��R�jշJQ�C���mݬ�܌5�l�h���V��Y�����+d7!�+�ytcg٥�ɥ$��㵅{���f�����
D�Yk�/�S��S� ��Y:|h�|X�K�5_�M�h!���0�I���Eޮf��� ]�q;�u��c��FGŪi��l:���~�����]�]�s�=���(#n��Q��")A��(5$�JPm��(B����fg�i���"���/9X��<ရ\?Ⲋ��/��ǋsӇ�ph����$v�[SG�O�̅j��l���u��J,�^�L�6�� =���c��Rߑ[p��z|��߻�|��~K${�g�?�:��l����h�H�y )~��Uj.nǥO&jqꉔ�j�#z
g1.O����<�I�o�������J��>��]�%k��AW뀀%֦G�'Qgw�S{�����q+������<41\��Nn�BW�[^&�X�pG�Q|**|�lk�ҶB�nq�R�=/,��qGM�RO�CK��8���L��7��&���lt6��ζ}������w�����Dz�\cҟ?��g��vߘ��޺��:U�cP��:�"��r��~t�H%�P�.�|VOK�bJ3�-��EN/��L�T����,�qo�0d���b��-F���;�"�����ӳ�0��7�I4���b�U�Յ�%V���-=�:�/Q��x2�,!5��d�/1Sqd�D���z��dPN�6�/	'�d�bg;�OUTRxk��d�ñ4�ݷ�A�R�22��� '7]��?R�}q��`�|�H&"il�[�k������B
��h����B��Y�l�p'�CZ1�Nn���7��w���d͟M��A�����,����'ߌ��6�`|�h�^n�d�ǻ߾��^CdZ;R�f(�q�Oha�̓��M)<�4�v`vC�g-ֻ}��ﻓ�b���QJ'H�GC���(�\��	�G��$h;���]��X�G�W��*'l�_ [m�Z�D��h���4J���PK� ~3R�
tV���6O󌾶���j���CZ��y#�7/�r�)��p 7���[�yEB������e]+{Q������|OJ&�B ��٫W��<�~�L�]�l�0�uq7?�S�S0��2.�z���O؂��aaԐ�H'8c��������ޑ�&*nLΦ�g�OZ��^���J,�S+g:t����H�'u5,��'w舷P�cD4\ݼ]�S5�ҐSz��;���1kF��s��/L`�� ��ݪ<�-�G%h���=u����;�%�������+���7���7z��S�|�~V>aƾ:P}E�J�ə-1�I�z�=�*S����`����3����*P$�D9�\~���ܜge{�������"��xI)'���3��}`v��V����mU�����,Z��hWJ6��)T)�<�N���4��b�"�,E- ��;�d!C1�������y
�"!�����)���&��7�S�� �(�J��\��*�?<PS�>.O�;Y�#&Jv#n�VX�lw��?�,�x�/�k0��|>x�3O��X	M�y����Qm��a<I��mZ#2�ngw���=���?ٲ��	�=�O@ȢH�hv5��`�q~�\]]���u�^&�"""bze[��!�Z��T��X[z'\���~���ׯ��=�u- ���Y��_���lDٻ���p��2|������'�(y� QP)��^+�g������&���o��8�ǾD�c�{$[>�/�j�Yh2n���̠@BY�s��TZ�m���' �<%οW(�>������#t��p�sɿ/�m���-\)CΎ�B��:��x��E�f)g�+ƳN�P;������Lt�2�31��e}?1�����Y@B�S��;Ap�@�;&���1��g�=aL���[���F"sx�?[p�1*�7H�H�$�PF1c�II��KW�n8z@��"9� ��^DQ�?�	�i�%tk�lte�Ir�ݢHaO=F�ac���{ɟ�VPQ�0T��"��Ճ&wd�cu�X$��Im��ΉS�n���q8��1@����Zi�wG^:έ���$<y<������"�P3�_�]�Rd]�U�I)w�|]�Q���lB�6��I���|�Ģt���a�.i�o)��w�p�Y�Q����SL~�<�#Lh!���s�0̦r�De{;�@�6d-�5Zya��Ӯ���:]#v	�;E}L�X��)Қˆ0��%�Q�)��~�GC�������%gM�5E�[�}
��W�S>�{�1ո+nx��i��>�K�
�J������.~���g����-/����Ơ0�_3��U�]�l<�?Z)�j򁻋qT�V����1�A��5��i���v�w0N[����R��x6�x/@"�/��6�M>�3�|��*���My�V��*%�4$�g;���^��Ӹj_E�V��			�� (�C-<�0�#5��X�V�X�^�����q�{8L[<�N����W�^�(�6�<��9��6�H�o��a���w$��M�=�y��Ag��v4�Z�]�x��s��bT\p���[�=s�$���O'G1�)TN�tZ�m��U1�z�4ǒ�\��v��]���[��mCA�����("�m��(��"Z�;�.��{|�.\n����CW�;�j@��#ֻH|�����N�<�o������Z����\L�w2�����gP�M?�[l����>]X��Ƿ��t�P��:��y�\���v~�f�vb9F3�c�sP>F�<�ٯ{�9��OB��.ͯ<#Ge��GK��U�6o�X�?g�dV=��Q�߻OEɗ���h�Ѣ��:�C;	2Ol��F���.JJ�q�n�7I%�h��1c��iGU����m_��Hʜ�wC���O��뾁G鿾���5�����i݁�p�ڠ��H�zEg�W�[��\t�bcB'n*{��^x�*V���p~�g=D.�h�·%'s��n��}SS�nl����!�m�6�9��8Rz�4����I	c䥠��h�����[�KU��0��.A��4"ZFX��>�CW��6�(`Wh�v'�"WL��XH����~���M�<�'�z�<��L';C���^�����qz��Ҟ;����e<���S�xv�b�8�K�e%U��B.^��iy)wr��I�iў��da����O1�N6#G�����N����u'�ؕ�Q�?�I��l�%�v73Kcҏ�����~jX�&_дk�?�_] ��W0�m��K-T�Ë���
dE:���,��*�1�t����Q�^j��|�_����D6���o�agwq���RQ�ź��X��n�ezm�.�C�1p5���<���5}��pJԠ!��T˛=ش��
���K��Fbsr�*�Ì )�n�
�\c-���A�֨�$���'����@tUp��2*ȏS�m��BT�}`��(b��xAs�;(��;��uk���O���%kԿV�I��w�*���I���]M���L��3M�k����)���=�0� ?�(�C�U��I����ֶ���;}z
�P�V�˳*��6)��5	2�W2�P�ݔ�2��7�&��������YOt�Ms9��C�H�7'm��!�Q�����������Hh��g���L�(u���YG�b����;Ȫ�,Ɗ�i���ס9�a����D3�4���^5i��ަ.�L��@���_Y���i+g���U��_��J/��}B~���֊�@� �g�J����U���Un*��¸\5��p�lH��w*jsq�!�8FDU�D#��ʶ�B�-,���bI�'��X�#��s2�IC�|����Z���&��%f�܌?"~a0����'!.��J�(�����]Zv���ȇ��ts����k}~�ÇF�5�W�$��G�}�/w�ҊZX�Mw��P���o6��{�Tq���Ӧ����ܮ����3�"@���N��]\毾�2*TGR����f(!y��;P5G<:Cƙ�K�$�A�?*CnҲ�ԭ�;+�'��]������β�bS��.�\�|��<�l@G�o�T �	X9)�Hߏ�Χv��O���r>'�Aְ�i��cp7+�������&"�`0����*?��;��X���~R�U�I�~&�.������!ߤ
�^6�����Oy��/��'o>!.�-�D�9�һ�����8���4�	.Տ/����g��{����G���Ҷ>�ӔN��ׯ�+��9EYRqS`L�El�?hkZ�t�p5�Z���$-���Dq�ݛ(eX[� �YfX�vFg��q�f���X��	��aawqE���'�+��P�nT�k�8p(�/z-��e��oyU����W	\�����9b�P2bus�R|� �}�˄>͌��p���G�\�2N�c���/8��9[Fq$K��XZ7U�-Х�3�L�Y�0"cx6d'��j�̞���u�<^��>�*���@*
�~�׺XB�R?M�腡�S~;��RhO娂?B�blo��%%��t�~����餕��i��S�"�	�]v.��"�w��^�Gs4�	��~5Ճmë��C�uy�� �����?k);e�������)c������(\���TZ�K5�����W~���&��N��8���q���W-O�)�^V/���3A;�M��5��#,z��*�?E^��,�N��) ��[A�4P��f�(Ai��䯅��P<_�Rhb�R��j����+�ߙ�׸ڍ�<b�\����U�����y��I��[~Lr�����Q*V��N�g ��3ݹTS��{��O~�P����OQI���p:��K�i�I���ic�b��4���q��5�:��:|p�v�����@�Z="��5�&�3`�!�<"X��]J������$ (�"=�w_��(�#&yu� ����h�Y-~c�\����^b�q	�R=!J����p���ջ�T�%�v_� ��7^���7��{F������Ld�`�o`��kl��p2%��vLE�9Z�A����LFDG¦�>���mq�{#s)i�DP9+��d�����G�l���i�2���&`�
��Cư��m����'��G!��֏^�L��|���R�J�<}XY�^�j�1�¤g0����X���ϋr�����ҡ���Zjy5�t"��.�r`P�15|!���9�𻆙FF}@t��V��^z{��fW�ۜbKD�O��,�߇��K���;�y��u�-�k�����D`'<�%@���.e]xz}��f`9g��2:W��Oc��s�]\'������Y/Tv5��o.!��F��ܤ(!-q��ܳ\����%ꛊ��p��̫�h[�/�uMi���v�5L��Ŷ�l�=� ���;d�G*�$5�}�[�픨��^�9a���	��y�n06�O��5�����bN����*�^
zrY�Q.�,�ۘbQn��
P��b�\��4A�2/�%�J�.��^S��Mvj$�zS�M*�B��fՌ\A-=�9��K�W^B#7F�~���[G��� ��^�����̓v'���>�6J�|���Bsu�_����XQ�❍��!*�^������2�B|�$"R����FM����~u%W�g4G2��,/����:�8yu��ۊΚ���IyA�^��u�$�U=�Z�ɩj���S�B��(d2��
sD��R�e���A=��[8䢙�5py��k�t�9!G�H��9V�nʀ+���<���\r{�c�'i�	�50�j�Lx��ԋ�$|>#�T����+
�����~�Dx�L�B���1*zb>���(������^���~Z��D��������(:�~�Cn���$}�=iXg�WF	1�T�Ű6��"v�~fo�6z_�'XY$�S���,���ʾ�1�D��i4�����yD��J�ly�4��%�-U�p�����+�[���p�����d�$Pn�[���PLŐ��_���`םN�,V��#�3�Rw����L�!^�<u�)�/�h�Oo<��`ųR(�ӡ`��8��F�_�O�w�o9�!ׯ��� 9��lP�������T>����4�۶��.p�O�tZ�]��s��dOGP�c���g(�����35�V��>x��K����ǰu9�����0���%l���K� H!���TP��p���:�]v� 8��$
� �!�����g׀�� �0�@�zg����Ǟ@�)����z��14�ґV�S��>�VV�+'����?#[Zp(��V������=��I 6�TثF��T!Y����"�9�L�f'yhnVN����p��m��7��lx��1u�/�ьe\�̾��ǆ�:�p��l�����1���iV�p��h$�Z��T�B4��=�.^�Q���R��n	���FKw���yU�J[W���1j��Ž�e`3V����'���)(��^��i����r��9XMMM��o	����(�"��/��$GL�+��Q�6���jj�7g0i��m͡!�^x!/[{Y��/L��(|V�N�}�'�FLR#zP=�D4�����V�o�Fv&a!��St��89Y銯YM�*--�v����*�Q�._L�!F�+`-�e�C\1����J[f�j(��̺o�,ԩ���NP��N,�����քq�E�1Ο��?	�SƻYr���/N��í�/*".��8lC"����7#W��q�4�!e�K���1���+X�'o�CQ4G�E�SN%/|}���-�)��_��&�s��e����O�� {n��1xC*-�CS�ͻ⢊��;s`�$�G>
ӏ��.N;�sP�V<-R����b҇��$�=��V={�0��d;�f_:9�3�$u9m̓�B�ܤm����_P�n�-��_��~e�ovʨ��U�(�C7��U�ߚ[��/�|t�`#ds��H�h��t�C�%�nD!68�CV"��m�C�KJ,���J���S��l�*9��SC��7C�nR�⴪�٤��u �>�/¸�۟�/OD� �ߨ�I���ͷ�Z�j�=��� �Թ-䬷B����7��Q�`{_��w��\���^��@p&��p���e����������I�x���-�@��x/ہK�㖃T���~1��)J���?���;�<�amd�:�5�@�\�T)��jU?u��8��� .�#�y��}�O���{RULAW�����
k�%H�����d�8k�������W
�ŝx�F�k�8Ĺ`�S��&�F��*�ɐ*��_�E�r�W���-#@[M�N�-� ���B��;6]"  �y�՚��F_z���Ig�������u	�������vR�Gj
�c�9�`��k�	���LY���r,D���Ku�ֳ(�Iı�0 ���y����r�͟'���bX�w~��t�-�~�T3�h<X����P���f³�� |� ��E9�C�dk�\թ�����a\7�6JgѱJ��سȤ��D�c\�_����<bM��kT�,�?\����Z��W�J� ^�p�JaP�5����+��3.��'��Z2?�<k�p�����b�f	��j�:k����?�~�6��Ȉ��/����G�F	�Y[�'�э�t���)X� �)��_O�����wM�����L {m�g�r�)M���sa�jKk�T�HE�%��׾��ݝn#Pn#���*��bZK/���G�s7;��X��	����G 3��W�'�����;]+����諔ߍ��X�f��4p���l��*�Nx�S,FSkt�+��C����/���|L��1급"wKv+4�KYͽi���>���ve�p>�X��:,��S2�V����D<���B&O���e�䃃��\��Ӫ`���6�n��$��v��v�Ϟ�;}�a�$m������������K�����.�~��Z�N�F�v��棊��F�����L`g4�ۑ�
s)�Z�%�2QY,e��j4�IkJ��o+_!B��%�G[�� m̳��h�������	�b^�8Kkي����<\����a�3��3O7��FN�/�1W������>�c�<��{���z�����q��G���~��%ʰ��|�21"ɉ����s��d趨:q��P���dw/^�D(��n��g�o,V7��W�\�]R��5f���6%�D&�^�!V�;8C�r�r�?Jy뱉B�F^�ie�'��غ����SL�y��jp��öao/w.�՘����*0�4ǧO�y�<M<ߦ��R�o���~��@3��Ւ(a��R,9�gB4�n��yU�q�h:w�gh��I@���R�~I��q�o[��%�rP�s�@���v�G�M����eۖ��-I\P�j��l�W�+oC����(�HYu錳��A,��0��E	<�/&g�t�7����]$=�bsnwiXֿ��������a����e�az��>Z�AA�J+�m&�cY�z�Ғ!1� ��\_@���^h�Ĵd�Q]3O]6r�G���:6
ߘ^1,jH�	�p���y�m(i ��w��P��;LA�7J�bm�����;����V����E��xBn~^��<T�ߺս4�p�x����Sݜ��Mqq}��x��I�����{����� ��5�|���ɭ�/Ռv�s7�s�U�)���+x�h�}"��X����9��ө�~�ڢ�jkH���;���M�	#��G5(�4Z�p�&�w5z�p`3����n�m[��x_�~�9O�V[J+�����cZ6�]V.ʘ}[u�3��2/}O�B�Ot6��cv<���GA�|�$6`ύ�r˻�k0�6�h��,C��K�7�ٻ���ؤ/�a�k_�cg�(_����3���j;�l�z����4%�4'y�F����L�I��_,��O� �:B��uh�xǌ�a�ܠN��|6����]�ݩv��S��G�n$r#�r�;�2��m���:�JKO���d��ݞF$�o'}��$1(Y����^��%�o�y��?ŉ��ߗnV�	��bE�;:S50Uxj�7-�Lh"�~F�ױU��[d����h]���G�����c��`��0�8��ײBv���J)�QvV_9\9v��ʗ�A��/��~'�*�*��G�aW�P�@j"�/#�"�{���]�������I��}M,�@ڢM��X�7oHUzw!C�pV�UJ
"�
�*'N����k� r��i3���%��n�L�c�%}��-�6���?tnO��Oh����m�O&ـ�v��$K�hZ&��z�pEO8X=��ޡ�GM�b�Hg��X���OZK�r �j�Ҙ�4^�kQg�A��x{|�z�9Z�������	G��m5Qw�B�$�<�L~�zA;�.�?��8�N�//88������w#�b�z���:/�v[��A^`�;�6uo�&���#tԠd�x�����Da���!���®_1mY�Ɂ4�͆s�1ڪ��S�/hB�=�6N�:S7��j'��RXX��D�{���J�eX�"����x)[l��Xv0�$*��o���8.j[]�ш=�����C�jW�j�(Bղޢ'��$�;T��+�z�1��$��h���F�ڛk����;�;��kK,`���"X|Kdp|A��Co�\��姚%�{q�ۧ��I_�f�2j�6W@��'ؖ������xE��6b�̘�G�]�)���D6���1N<\�U$9[��Tks�i�F���7����ģ����q�|��)����0��mÁ28V�Br�e-��Q ;����|@IP*z�>qM�N����O"�OSg)PR�;�5������"]b��I.d�����KR ��ab��1��ܩ/>�����j���S�lXTZ**v��c�C���|�z��pΥQIKt���Fy^�0�߲Qc�fT��},c�R������a�놇��T1�
��_Ъ���$"X�Na�p������Ru�9�K9mG�^oJ�u}>��v~^���4������K.�	y����a����B^7wi]*Pl�L�>�٪�.�D&t 6MG9�#������uG~6T��=��k'�T����o=���oC1�k��N�TC<{mfÄjrK�C��>�:o�"��mVQ���Z����*�]��rd�Z���\j,�csLZ�x{&�Z���p�:��xP�h�ݻ�uQ1�fGX�Q �x'o�
Q���L��S�5�d�#�GN����j)s�Z
~m�y�̖�����t�0�;ZQS���b��>��x�z�*-|��R�h1K�-I�Y���H�j>�*��/�SHk?@��r�F�g�	�W�Ge�#�lq8�- 2&�z��bR�0 ^j�(�*���2�]�\�����`c��
�|�Z�(ұgS�Q���h��pn��_��6 `���e��	<��ɒH'݊ŋNx�R�u��/k�;z�G���r��]9�G��?*��	L1	�8E��_�C�C����<�i?���fK'�o���?"���9���/XA��3�-,�HO>�̘�㌂P��#�um�e	��
Q���>�}��߶*��0~3����:�҅�׏\z�˼�`����M{�\�7�`X�G
+��p���a�;fp�!FPC$���WSH��>S���Ɛ���>�J@��_�6 ��UQ�m3���LK �*d�����ו+�@�U�l'HH.�s��̔M</+�OZ�,���6Y�}T`b�`������6�g7���AOfcå�&~���#�b�'^��������濝����5q�j���?M%�ھ5{`��FBAٰ���-�{j�R�����=��3;�"`nZ���K �밑v^ǟ����	�k�vVӑFgdӢ��Y5ݯ��$��$��q)�y�m��,.X<є�.�M���������k��	�M�qi_�:ۜ������s��Ś�(��(�@�3�OP�ET���c)��#��>�1�/n����*�?�,>���R��XJ�~?���0��qM�q�I�p4H�42RAAA��Q�0R�A�AJJ���9R�F�����y^�����s���_{a���i[K�0��B��P���Z�,��@M�s���5	_��cXǌ��j��o{�{� ��x�-'�s]�sv6�/]���ܸ���&�)��䌟l�bkРt̖b�t�G�X�
�50�4��k ~��$�6J���/g�I��3�����=c�Z������l3������]͇JQ@��I����%�ά:�~*L����U�"���A�F�8�W����*�K;?,�ˊ�%����R�ݏ�ؗ3~U�t�+�Y���}q���X]c��YdB�*-0�֢	���: j,{W+�S[�?��uM�C���`�Wo�(Ұ�I��`V7s���x�q;�WVJ�Ў����F'���7!8~g�u��!$��*��RLTA�c����ߣ�]^Ɣ�l?i���isp>d�Q_�_�0�C�wO2����$��3�Z�o��C�*:�Uͣ!�p�D'���t���5����M�7�j���Ab�'C�z�b���6�6k��g�U���NO�a�����*ς�ϒ���PR/���o����6�n�h���Qj�%/�8���l �6I�ԏ�W����#�|cG�7���g���_�)�CYg%Y��i3�jȍ�s�N��3�����J%	���u��B�.Fj���(���
������|�yM��غ=i^�6���@��T&��9 �jZe����"���g)�Oc���¿��tF8U��V_�c��0��y��5��g�F_��7`Et�׶��I���1��G�Agx�-��g�zZ���	��P�k3��玷V����Ϸ��x��!�,��S�c�Ƭ�R��(���Sp���H`*�>�qږ���&aEH�8�+��H�%�JYg�Ivu��L\���y(�o-����<{�$�-���1�&/�$|	(5��޹��s��ɺ�j39cā�M�g��ś:�:Ҳc�F���*1'��^M��=E��E���q��`�*���#��Z#�,o�_S����)q���K�]%�U�Ok�5)7|;:�Ď*PZ�B�V���2߲\�c�����uL�A��#|F�ό%�؟�K8���)Cm�^Z�R[*@��z])���n���}-�>y�!;��ĳ�}7�f;����w��4�PK)&��5����*~K��JmM�2.�$�>.�}��\[΄��&7	�a5��{F�Dc���²D~�1�C!�࿔� h$o�L�T����%�p������0�ܚ��:�:}u�!�n���L�
��/-��xIo��'�6+^5N��b�{���UL�h�(���,�QB&P�T.?�0kC҆�d���EzH�oM�5���~]##S�����x��pۓ/�	��7ٜڜ���Nm��/yB�M������r�2Z}W�,TJ�u�©�D�f���K�$i�+�m���?EUO��ĭ��}j�i�*�g7��݅�|����x�5�՗qR�\g]6[�29O݅�v�<���>�ߕ���M���k�Z虁�2�s�|,5t�w�)o�T�T*r�mG
n��۾��A� �>�}�MF��
b���q��v�R�y�G���8����zN��jP�aa:��<�]�K�5wB���A=)4�'�%�WN]��׌ct	I	Λ;]�j$TT{�Ӗ�e�H��[b�"Z��lu2��yNmկ���0��9r��Rp@]��ll��s�����Cm�1R����1&�HbwK?�í��W�Y��p�Y��$���T ���hۦmm�V�8E2���)�q��3#���~xk`{b��r���P�ۼW٨�HL�3}��rR��m6&Kbl���0�թ�p��wֹ��y��߲��F�ͻV�x���7�����
�5*��]@�SR����8=�4�}�$���3���l����*o�sx��Yź�LV����R-�K�=�Pk��^�UC��\R#�=��$�_���q��Y'M:���%�g��|����O۠�����%��I;_��vЖ&�S`$X�1;�W�`�L�?����l���K��zh��S�)'�ck����dKo���kG龥�B��a���4��e�*�\b��0��EN^��/r�IZ�-q6�i����ȼ	c\�=w0��N��q��G8% �}8~��-�g�a�
sˍ���J�(���3u���.:W.�|�Â��d<tMa�gTx��N3L��ǝE��	����I��MŸL������b�l����5����뺗���^�3�S�^�-a�(��Aa;Q�r[�
���)�˚�����a_��	�i��Ӝ(��+��A��J0g�`��X�h��6�[+
���O����"��G,j�*e��L7q�UR�E�HI��5���&�)��QzZ��l�Mq���|�sK��_��4�)"���$9��u�Au��
'�;�rܠfj��Gr�?����]��U}�]�*� ��l磈���\��ҿY�?��P��/ͺc�+���+Xf b�l_�P\J�O�U�e�UӴ�x��c*�7��)W� ����tO��,�� ��MY���#���i�+��++dm�����ѽ������Z��a=#^%i�j��g)��v����,|5���0����V(��p�7l	�6�Z޿�x߀�E��ƿ��*�C�o�q9�R��`�'�����+���x�ka���[WvN���3y�Lޛo*4A~E�s��q�g���*Rk*��C�`X����*?kd	������s{w�'��+�ӍC�TH��+U��\��s���*��A��p_�1��㬽����SU�-r銍g`D��ՙ��p�Tx�3��0e��[�����R�|V��%��ƍQ)���<�Q�:'�/�8��MEnKG�j5���A�(2Lh�4Y�X|�.)[?�ߟ	�,̌Q�N���u��@%h�H��5!|�e7q8\
��-;�%���ޔo�������]G� ��;���Om���QI(����c��a���GRUK�z�1L���_��L��M%�[�މ�O�3��}����d!L�p���6��/\�%塙L%�ڣ�i6��L���E��[�,?��8v/�R��=ݔ4��_�jd'6a����_�iT',''�5��5^8ED�#�t��"��9�u�]�^GUUL�}gO��&�N� 7;92��?�Z~0,mv5��72_�e?�Y�.BE�E�p\�]���iX��->���:S��fM�`}"%{PoOk~��e�U`u�ű=2=�U*P9`W�ct�z<��"}�i*Z�N�����\����由n��5�7y-���!��3��
i'oɬn=�΄7z�R���6��!�&?�lzMد�F=qie�ntɿ�2E?I��y����69̼�I/���ȝfMh���`�J�g�+��"ȳ�o@����i�?u����]T+���"��s�̐M�:!<1#�'.�s��C� �v��k����ѴE������֚� kڗ�7q7�X�����J�,��TL:lU� w*7%'+�集ć@��%9kgx-IJ��w;;�TZ��CnͼZ{��`������Ak�5^t�����R�����W��aW�06��3�φV	+���T�YC���J�,&;��|&�Jh��oĵ����äȤ�6��W�1
6��z����6�D8׻���~�7�Pr��$����<�L5�Z�M�k��>��cZo���*�J��;S��-����߉x��\����&�>��-��b?9~?՛|�������r5����� v��Z�s�q��˼X�P�?N�a�3����d\��A�+�̡���� y)
'�͒0&��O�LP��9� }��Cb�U�$�C�J
�r6��4�����7Y���,�u�^<�'�n-\����������O�HD^�&������@Uo�查���`�i,��e�Bj���g�tfmZ�f:��}!zbiG�_{^��V�أDĿ�:ZW��ӫ�'}��1����m��kx{W?Ȯb��03���sRs[�M���"�(�Ǻ�O���0-
���w�2��j�j_G J�����*P��Ҧ�}�NN�׻�'�1h͔��?��6��ӯ3�g��a���:���r���dra�J�
"ll�߫�>7�0��6�ɮ��GCKk �"����s��IO�)�9Qf�7e$yQ��x�<�3G��R��-h�C6UZ?q�y���~J���쐓(�1��z��㪧\N��h���Vb�(���e�$2�=�5Cˠ� �l�����j���b����a-^3f6Q�|�/�=�
n�n[>#�����:ӺW�'�q�;*E��f;�����Hmj�[�.3� B�ŝ�&9e���]К�D_��(��t�!� �A�o���۽c�b$�~����f��N�/�X��~r�=*0SF�����l~V�щm�inpoָɐ��T�9�q��3��>>����c�;$��	��\!���fFƁls�J�Z�& 8�P�ڗ������5l��~t�-��T����\�Wzd�R���RN�n&���%��U�W�wt�#&�D1!>�?��8=M���GN��nWh�K��b�Ơya{%�%z*v�K�M�8� z��U���L/�?����N=i(�OZ}�b!����`���<L?��О���լ;�L�!\J��/P�V�����ظ6�x�Q��D�ۧ-H&�M�ƙϘH+�iJ�(��5|�c�9�u/�ٰ�-V� �J��_����r{\�"n�'ߘm�P�r��}�D���?�8[���A�(i߹\��N{��ƌo�-�&�W;�ђ���{�vbR�&��犮R�3q�9F_!ҿs&�o�e�(�V����%�Ȍ:<$Π�	��K�[�,q|�y��LOw�2��v3o��`���:J�Ÿ2���` ��,�]m{L�����]�vOļVe���늕N��v���2d7uI�)��8���0���Q57������4˺&��u�;>�w b��V�4��I�;�lf�v^�!��n�0�0�@�����,)�Xb:�N�>h�����o'���v=b!3� �4�d�C�$>qvP+l���<c�W��Bj��֊��\ƅ�=�����R�+>�-���Z""/��Sd� m�<_��T���r��)��{��",��5��3�̬�S�"n)�04�ӧ�n��ejfC�]�Qw��p��w�0:w�i$����=� *�7������ǌ<9���@VO4�쯪����ͱ�����3\nҚ��bR�UNQ3��x?��0���F�^(+�P�������J,�"��/ �����������F/Ud�$��σ
��u?�뱉��k]�\`te����)����9ۄ$:6H�v��y����=]}�/1�{��[�G���0'K�A�s��>t{�Qo�n��t�M�Nf0y�l���~/�[Q1'%QprvBe� �C��hqՒ:�I|��)�B�}��T�)��ja�r� 5���o���53�6^����klkzٯ��Ь��:\�
*ՕP
�yoC�]Ra߿�1��~Ur@�z�|��w�%�wƟ��p�d��	��j�ߣk�-ß���Zk����l�����R/-H��W�*au�ӭimEMq`D:|���Q-k�c�:Q�蘇�ī����9��GK�a���0{T�K�-�)J�3-�5�Z5x��G���e�,<�7�@˳�����D�9c�~l=fܱ���{�
�?
�*j��2}���z�[N�ʥ�9e�%��a�����a[A5��O:l��t4,'U��G"���ÛYA-��+g���S�饾`B*���w�~��n6�y���_�L�����;�������T�`=,>�9�\|U��2}���U����^6�I�-Pfm�,���W�����#��!��������W��i!��=�J;�V�G�@������b�1�M��7t��#{;^���Eg ��I$9�M���/���zJ�౻��>2k��r��ُ��R^���L��i=�И�w����x��b&���ŷ y�s9׎��6�W+�=�����2Z�k�T%?EI��>�|�����ǌl]���B|��2$�����A�o�Ɖ���pU	A <���	��^�����x�.�K%v��%/�O��fr�B���>�|tx,�/��Œz�I�&��W��F�=�ծ�F�]�*k��i�_�6�������< �Hj)��&Ɋ�N�/��	�.1E^^�����0���j���9q�S�����V*��I�_����l�ك��(x��įa*X {����Wi�V������x��@Zӕ59��d�u�;(5��iJ�*�Qs�-��$9y+];N3l�����}�[�8�$���֚Pk�I�/h�Ǌk�2s.ˮ8{��il�c޷ϔ��W�y/��um#���#�Q����"<�#�~�y��d�)�f����j�	
>���eabs�׺�6��>��<y[��������,�i��<[�l]�m� �J�����^�#�S�n��*���W�q��B+f�S��3+�C���KmTJ��3���T��h�����z:�o�҈뎞����}��$�4���/ 1�n2)�m���0�\N���tM�y@�g�8'ƵMf�m�l��r����ĉ^+	l�)t����Dv̥E����R׶�%t��XYZ� P]���z��ɩp�S�ɻY��1�X�+B��E��u�o*�Z�*��}���@�<�o�V"��M�&⌇y��	O�~�A	M�Ҵ�2�l]� ?�2�B�Zc�Ŀt��*<�Nko<-y:�r�2꟤[��{�)���Y�D$�`T���v*�]8�#w�O��@BDfm(߈�噫b��HYT@ʰ�%Ve��$��c%�}�&���wx#�*y5�3u�>�L�eYo�M���0@|;PK�,�I�7V�"#����lp�b��2$�����d�P*��תojh"̥�Jd�锄n��Oq=�O�b��ӱ(�Q3���޵HO���Sb��)�
P�tO�; �JEy���}�m���Gr�su'�\	�t5g밣�{x9�fHD�r�[�rrkJ����};��94N=�?)3=�\���9UN���	�տmˬ�h�sc!�.)&5�f�郠�姢����jS=O|c!Q?��?p��+�6a�O�p�QS��_P�З�7h~(�y�D���` A�t	ܲ!��]G3�P(7����Y�pF��wc=a�iX��JG�c��|��|S1n��,UjO��B��`�w,b�r��yRo~�aVk��U��-��3��G���<�1-��E��������'�����Y�Wiĳ,�5??��A���/���g�)�9"��(n��)�˗�������JFF�_ �x(�p	�I�x:�LՏm��=�L*A�X^g�:��^����ۀ^��>WP�e�Q����T����Tf��cp��pQjq�3#J�ŷ�����Ax���ui�k��^SVr����|ɂ�5a�Ȁ��w�6�K@&�-i�뮣yy�u���ó℺c�h.��	��'���<��s%�s����a��ɤ>D�\߮�8͘��c�;�yh�gj�&]��O��A�7��m��>�ҿ����egg��ܪ�|����+tg�I�a�?����ԫm��bI�v=#�jf�d0_W��[Ї��ʬϞ��0�W?h!�N�9�$�YƲ�o�L�+���IF1"8�bޠDo���v�o��MA��@�
L�>s�E O��1��W�����bk5r�>2��c��\Ƌ���=��:m�e�n�R����5�k��r�7$k���醕�t!������r13��(����v�z�Є��9��=���Iċ�ByV�V�?��{EP�-�5󛊸�@�/��U��v�����ѳ.��D��k���~X��[j�>[*_��go�e	fp�l�'��	A�0pGUHk[�91IV��S��S�$҃TZ��dg��	���ȺR�i����軞������=��G�ko{��Jż��b�eH���'����?�� '�v���܏�+?������,dg_�mM��d�������r�]W��y���Cʪ�ʾ)�z�� {<iբmԿ�)��c��Y諪u�$���f%흟%�g�d��ax�?�8W�W{�O���(-"�0W+�j�������S��BC�7���-чݙ,��U����Z�Ϻi�J�WcW��=ok���U[?0bJ��7�h+�G5}�zSK0��a���V�z�������/�/f���h�mI�)	fI�E�\;�@��
s�B�dk�z�_U�>v���T)Z�j�0�߶���vBJ������@=bJƮ�ts8ʴ��GEJv�#~?��R��MJ���Rijk2W�cm�wޢҚ_�j�u�ĝ�SEǼHv������Nu^��q�8SsQ9���)�h3?�|�y�wt��c�.RC���y@'�����o������r{O&�t��R�M�˴���L�=�����1��-��R��*&pP�b`k�SM�i�XOU4Z�7M�S	e�������9l��U�43ad�]s(hW����L<ۼ@�aSh� ��M:wOX��M�U��v�:�c{r�y�5��j� ��9�ZU�TkB��y���9國ܢ?}B�(l�K)�����IĦ���*ٗ�ehw�I}_��i3�����~��5���RB��x����������]�y�C��Bbɷ���[�9�9=�=B�HL�^�^��1e<��p���Y�Wb?�c7��Ŭl�e2/�mߺz���p7x{���o9������$���5-�Xg�"#�>L�Z�]
;�".F���f��,�
?��K�i#��V<���Qx"�{�M�����/�m1[{az���#k0iP�S�āw�T��M^6�����l��'���c����� 2U5U4���S*�fA�>[�u���\� �|����^y���R�t��Κ���FQ1]�wC.>���d�и2)�ٸx�}�9��2��%=vo�ظ�S�U�2�G����eY��Y��@sf�^*���T�#�]�M��[�q�Ƚ��ͫ��k�"��Q:"�ދҧ��TE�5i�AM@A�>������������8,/�sb����R��Fz����8Qhi�i����A�&�� �Pg��DRu��;�����J�po!�j�vꞫʏ /|6�vݶ�!E��J�9nR�7/d�`�݈۠=�^7�Y�q^Ʊ�����S%`�ɆO�� ײ��+~�m�Qn�S
��a%��S��}�T�EJm�3�8}��|Q�aW@�l�����ܠ�q�_�l*��9�<8gѭ�){�#�"�0Z6 L���
�%�����Y|f_�[L�'��)�^�9=�J����a��	�Gx��۰q!�P�/���h��s�Sܸ}?y鿷�v��^�H��W���W��Jv#@�#��+��@}���g�ٞ����	�%��ê}U��[q�:��&@��PS�
�,��D%ˊ�:���˓����qW���ZT�$g�����d@�?|kk�!9��8+�/�:���٠�-���M1�=�Hzá������9dNl��Eq�*��:�ľ�������5t�h�O���ܜ����4�$!�~��.�\�nkJ����	"���O�W�-?e�&r��O����\�t�~Z�����,932 -����켶� ��՜�K�@fjv���aTZ鼆���-6T���e*" 4?�2�!���$ K�N�k�����������4:!T���i�J�ϣ�j16hf����κ���T»|�gk�j�w��@��s��P�Ҽ�s5jYݱ��WљT�����}��>�|T5�TV��Q�-c�����:cBn����[�+q5�me��N����+	l����aʈ!!쉰����)�u_0�"�1�U"�BpU�j�������Z%�	�y��� Z=#�v��Ob[ͳ�( @���(��c3d�} -���?�2"� �<��8}��Y����$g�*Û)�6'��b��,�-��F��¦	z�|b���&�����U�a����
k�����m�T��ۓ�owwq�%�T�)
4,Lᾖ�r���
��T���J��k�c�b��!|o��qR�[�m $�������f>Q��ј|��$Q�J�&��S\�������yP�Q���g>P��.�Iq���ʞ	.�b&1o�N�l�ܼ��PV��Ӊc(CV��3��p �h�p@�ԣ���'s�?#�DkuH�2ȽQ��׺����U��������{���?���%�`����`;��(��:t߬b{�)Y���K�[�4��(�h
�lGME�OZyHx��\��fLet�5a���v����;�b���Ey��fu�]݀êS�ћ]��jh&�?�:I��y���Ϸɦ���./(���,@�3�,әz�0�v��ɉXd�^�ٸ��7����N�d��n��fR��{ey��x��#�dwU=F������eC�dt�����\_ �ɚ�拳�;ۉ�6�뎵,V�.�٩�T�Oe��VK��?�M{������iv8m�a\��n�]v�?ͦ���[���<,)ꩩW���n�ӷDüR�c���>h�H40�R �� �+�w���N�"7�x�K8]������V��t+q�}��S���;��`��%f^�M��������Xd�r��BX�:kc����Tڵ��;bϾ��?���z�=y���qKV��C��<L���b=�J�S_�b�C�~m�T�4;è�^�uvx��;W*�����mM$hA->�m����;�W�npF0��=�t���˲�4�n��T��>��f)J�����1���]�B���#MH�{��L��Et�#`�ά��;6�Cx6��ϙ���vqkU�$���guв��̞r��i �8>��F9���O� �[9nW��o�¡U4�ʀ���4�ۻ΄N���&4�/>��i���Q���b ʫ�Id��:m�\O�Q�̬ٻ��W�:n̡<Ǟs�niZx��$�ޭ��m�G����.=�daǾz�MOج�x~�Ҥ
Q@��4�K*Gi]�J$NJ"��0�FP��/��+}�w��K͚��)�pUe�aB��}e�7W�]ښ��5C���av��� l��!;|F��$u�ĸnv+aQ���>ݦ����N�vx>@�[���}�5�M�\]*H�A!�� B��@da��%�;���V6��>�f��h	b1�NX,��6� Y9��$|P�VT������y�����{�Z|�%<!��k��Q@��16�`Mc��g6R�W�Y�dnɎ��JVf��%�GqQ�h(�լ�w�^�C1y��ڑ쒉t��v?%n�̋�<�Ƣ��Q{�:��� ٝ�=}���-۽YU���c�O��$��u���'��c�৚8�m�?w\�miWt��l~M�S{c�W�+ Oi�Yw�(�R�j)�h�q�5�\Loa8��i��[��e�x�}�J�w[�r�a�U�L�r�a���ׂ�����ֽ��Y
 ����4�x�[��������(��me��y�/���D��a�@$�`$L5����_���'ӑ��Q��!ela��c� 8�Xn�X���Ӿ�+T�/41.�F���?6q�,e��#����-���%GT}��I�)���bI��M�Z��'�I�$�6n<x�L�PЛ�[w]���;�8�ӽÍW���>�P8�]z�ѧ�?x9P�V���i9�~�[@�|���[$� ���l�,i�]���AI,�J�	����L{V\��[�&?����p������Qƛ�e��o��t����M.��Q6�[x�-���@�KW�e�ܹ��3 �gޓ+P���OW$P�Ж��Y�Db~�Dǿ�K�
w���{$=��cl*5K	�����9�\cOy��vܷo*�irm,
�tdg�����B;���|��Y����A�Q��^�}�#Ȧ��"LV�O��n�}�	Բ;�Vm�ޓ/>�`��$��Ex�M=�[��+Kẇ��1;��縴E�M1��w/(�T�(�]�9S5(�c{l]Y��w�Od���tc4;�fV�k�"�ne��O!��*Uf;,+�<�?��W����۞����/��d+3�e�]a=/��yӺ!�3��o��^���KHS�L2�d�>�{5>iA����m��F�*�nI��_~O��;&��	ܬ�fU�U��nb���0_C�糒j�S�^Y��#9�''/&���}*Y*!��ŴBX�����~�D.;5�����4��D_o�rb�ݮ�!����<��m�=�{���I�O���l��S���H�������Ux��J��m㣋O ���_3�������n��I��,t�X���a#��n��X��H�zL�:.D{��eW�I�!{
5���ux��۫�/�~U�d���B	��C�xU��Z]"�g��!����M�"U�,TC���&��d������\]q���J���
T������-���?�FN�S�͔�=5�;��ZT�x���t�_�f�4�����ۨ׭��%<@�Z�+��9;�Ε���s#|�.W��,�:�|�o��.�nI ��0	
�(���;C��˃Ia�'�"���?��\*�h�ď�����ߝ�����������p�k���~��>7�F$��ҩ�۳n)A�&�H�u2���o�E�y�+����	��fo!ӆ�`|9+eWO�h�%����
�ﴷM$�q�k�7&�ohSj�r�4���(ekIBd��M=�42@���v�h@�����R�	�L��tND�sפ�E��Y�L�o�o<��R�<J�6��.=��wC�\-{�?�S�P욹媩��X���H�����|��n���n��җ�vq�{m+����34I±>1�+ɟ�b-O{��K�mha��'��@����o��T=��'������A��X� )43!�?%nϚ4� 0T�ļ7�D�"��®q�]��-��j&�z���R���3�P�aS�YЩ��^�D�զ)#�Gϓ�!;N��Z�2G��r>6�A|W�y��IQ���-�o�/��ny��[Jl�y�H��f�������P�B���!1Z&���'`fn+F��wA�� VV�<%l�:Ԥ����ٜ����A�����@
^\�8��c� �5�2��*6�<V�� -{s�z�Y$��#è�hLR��#�U'Z*U��.����K� �o�����3Uq��5A�����O�0+�I�2|>���;�ձ�3�y�}����A��ŦM�#)Ԃ����t������Ǝr��ޝ�"�> b�kQ]�NC�� ����ȱ"9=y��8���HuN�u/�Oj8}-�fS�V]0'��3��꼆�ӱ���9SQ]��e�s�gO`>тr�߿T:���G�3&��t+8�\{�O����Ck�>�2�ꐞswTW�����0$�0��M�)�9�p���h�}��噯p���f٫�[��@����SxC���V%���PS���a�X`p�D	F�af�#8nt�"��B}��Uy�I���d ��`^������2��Fa�BͣiUy\���w��2PU/^W��Ϫ���)x����Ҿ ���`T{�@��+C�,s>�<$�4�j֢�ѐ]�s{	C���oWl.%B�8Բ�*����l��b��{ܠ��f,�0?=���5��6�$r�n�F�o\˦ꊋBy��D�F�zk���?�P�VFi�!B	`�y�/��6wQD�p������β:(|��(�f�6���Mu0��.�{��p�n#�3e7��w�������:�T\=qڂ��t�E��s޹tb)c��W��8?���`1u�B]wz� ,��k�9<��3��'{z��ݕ�n�Q��Ϻy)ț��I�����!6rI����Kkujy{�[8��aNy#m����~�}	���0�e�5��H�������C.�fW�D���|^�k�o����� �V,��a����ɫyD�ew���"[�)'��g=��-�ϱ�n�)N�`[,<E�3-LC�}���F����ɨ�IC���T���;n�>=u�Z��wt*���I����gX�O�/7ި�N�=K�����H7���pտ8�}��5E�y�h��E�5���2�@�|�8��n)��x:5���-�������3Ц�mu[�~T��
�ލ���^$7n)����h�s��~�9�r`A����_�Cz&ϧ+4>��ֶ�Ks�oi�d:��k�ҶE&�<����=�B���{�Ő�]���G�,���܌�l?����� ܸ���­<<�Y�∧�Q�#�, U��V^��� �9v��-���{�O�#�Zg�;�����C��nK�(7k�{����K)�_�!"Z��G�T��%#�� 6�C������BiqG\�Dj�u����e�{kU�ƭ�An�}e�������9kYm?���\�E�1�Fb᤹#R��SZ��ѻr$w�Cg�A8�u/k� T�9��U�<�n�<=����'N�$�k�DZ�m���hn�aQO�g�We��@\���4���Ux�}Ĝ� �F�I��"a��u��ۃ{�l#@zF/I����^c�9~>v>��J�$�`$ֺxg�x;X�]����|�*
'EC��/��{)C� ����Rv���k���x#����_�=����[�;��*;�u�; Ⱥ�,�	J˱5�\�\��9�NV�3N�� ^<}�O��}��i��/	g����NF��W�$�A�/��^x�S�֍']b���X �5�i��+�]1��+��Ŷ��H|O��*����cSO���t2��O5�᦭g��v֋��![sq�}S�2ڽ�.��T�qֱ���cT��	�`�|���v��2�bf�����<$�*�ɠ��H٬#&�dq��C�bj��e3�N{�L���3�6�tc($��iB���Z��z�7]�^X����^E�6}zD�y���j��sMT*g���,���
���A�Da!zh͋�������&�xeT�"�8��Tȯߏ*`���f>`Z�(Jץ(Xr2x^�*�!�ڠ�j���j�C����vN9�������|~m���5���h3�v��%t:0��N^�b���W��P�7|�?��wL��� �����}C���o9�6)�urZ�r\n�DD�� 12 ��/=��ګ�w� �ۮ�
�y^���N�����fu�k�Id�ܼ-`ӂ��9��:�3�x�ͩ�i��$ز&���x-6_d�ߢ�N8/S8�k덏�*.h�G�_�flD�aXޮm�sn�n�Ӂߡ�>[�u.���;=�?���
6�t�������v��a�9?���#�	)r}-�U�䝂�]EP�ww�>��A�o��3��ǳ��J�4�0ΔYJ[ĽX�HYfiɠ]�`ga}�gܜ4V�9�?���d�༞���X'8K;3@V�%��:"�w޺�؆����)IZ��ݻ�պ��쎨�y�N�ȳ���>H+"&r��O�͙��e���{D4�a�5D�����lAˢ��z�Mڽ����;���B�?~ך������@K�+�}�](��~��w�<��7P��j�ok�8�Q����&.�>h�M��Sm^M��ȫ�Oϴ �GL��l�J5@�{/��#����ў���ǟ�oPKڇ_C�)R��0�+1��@ԍ��=�����/�f4�߸�2�b�m����=�	����7
�0���op�]Gj(Xݵ�^��4P
F�{�Z�+��p�']�����8J���!�j]��/��f�g�A�ݴ'}u6��>��R	�Y�������eҤ��뉞�k�b>�tcL� b��G���m���G�f˙�i��ꚯ?���6�6�zq����~�ڴ�e�kE\� �_`#�ųj�ܠ�긻3@�ӽ�v���X:���'�~��P����pQ���S#h�o�c8��	`�������䙏4�V�NKBF����2[B3����&�'��(*�܁�����w��i�H����07.�n��N�&��(��"�\i,�mj�*7�vOV^IF�u:����ȈC�~�=�0w�
��"/���^A�S#��0�Ï
�o'������ϧ�^c��<����[m��a �-��s.���=�VLa3�Ą�	P{]��Z&�wbuG;r=q�����4,���9�w��f�m��{<Rk&� ^U�P㮣2#�,���U�3�M��F���B;MF˚��}���]m]	=V9[�}���4�{k��*��O���V�ܿ*{���4�m�9#��Ye��K�A���)a���b%��I�<F���kƳ���)�W�u������-��j���P��ܵxKphq�
�(�w���Bqh�Hq� ��C�����}���+ɑ��̬Y��Ι�?��6�1�?�k,�]G=f��1�0� DI�7��u"IO��tBӦԚ��;�+�ߕ�oE��m��ݚgt:je�W��!��/;�h4ߢ�j�g��n��7���b<��ɑ�eş�I,�B�'�2G�������cp<���5�^h���� ��F�X�V�YE�Ѭj1o/2��p�6�d�~D:D��mX���+^;x?Ecr5H5�o>��ݢ^���|'n�h�=�Ck_�w�w�'�@t�o���"��_����PN�1z��*����D�m�s$�M���e^��yŴ�4���Ü׌�`��t�a"6� �`;+mS��8J��`�єM�J$YnA0��&R�۠�o�֓Y5�ni�0_,""�� ��}z���ē�@D�@lg��x,�.�Љ�m���VK$��f�Ǧ�Gͻ�pQ7���m�)��63fS�!3XK8]�ν�F1E���O�|$�B���Vw�}#�6^|�Y$Vd��Y"L�ǝ7���2��A�6�;��iu���� �e� ��h)��j���.���0��;n~��f�3���� �yӮg������X��Vb�5��N�W��g`t���˗��Y:A{j�/��\��NL�����c��-��+f� ��	Jv�,/-��hY���>b���!����T�C�q�+�;��|���
P�E�=||�e���x��}�1�]��>�	E>��	�E{�I4k�O������^޾������$�Ȅ�S��,#�Sz�Ƨd������>�����i�9���t#�Di'�KSE*\r��eA�}Ҟ7%����$:�����ن��S�t�g�i����S�[z������I{B�gg4�E4 ��y���]-،��SP�_&�n�dB�i�W�-�V�pb�����ŒX��2��+��]�DfVgz����B.@ct���6$�˙fI5�1%��⽘�?�[g�)�'���5�:��i������:����9�J�3�RUPJA�����L��_�`�6]Y]Q݈!b�÷8֦�ē�2B�y<%_8S�56��;�='��"�կ:�{.0��s\�3I,Py�
���g?���_QC0�$-F��	����W����-������c���ߨ��b�T��i@�Wu�*��~����(z�=6@��an>�1H�s�h|D@1�a��$�a6�<^��p9{qBc:�3�&R}n]����͇E}=�L���٘����T�Ң7'�Ct�}d�P������R��B/G�:�-��7-�S�M������Z,죩i�3�c��i�+V��Z�O��)K��:��1�.Ǐ�п�P,O�*��I3a⡝ʉ��w�"�}�*$]��+�L>�^��>�E̻��^^��^��x*x��Jh���cɒ}k�v4T~�x�]�d� X��������H_�Q�Eϲ�o5 ��f�u.�e�r
�
̾M���M�Q�;�v�2/��`'"�
�Mv�;v�#�-��?����cSl�pZb-Z���Y��B�Ζy�BjN˂�b*>e����\:�\ �W�c��FŒŰ@�A�٫�[��P���y�[�c<5�(���wHâW�y�Ns��$�5˂ت
ii��'�,Y��<�{�6�d�U%��V(���  �)�����=\� x�=�UB| ��L��׆��"�A@ t�3ϲ��r�e%��EQ��z�$��M��l�}��A�S�f>�ʦo��p6-2kp�7�s��i�����+�k���O���(�5��5�s���Éi?��ҙ^���Ȍ�댾Ǔ�?��m�y]j&�#x�ʠ�\�C���l����4[ S'd������x��u��y�K0M}�W�
��ON!��˼�����7r_���K��G˷��(6�p,U
�ү�&ė�"��5��W��  6{V�x���ݳn�U��K����?b����@��\ �)���*l��f�xQ�l�q����Zj����Gbh�I:bZ����S�N�Я�1�/�!�=��^h��Ӳ]S�%�O��\�o��>w�Nw�c\�;L�L��ed��
��.��̋���X��* ���o��>���V��������<(�B�8H��!���[��P{��cP��.:�� ���|%t
��v����ӏo��:���M�����̓��+o����;�m��t퐛d�e��݋��KE���bA����1�\�i��+��|,��c�jwsci�N?=��Q�����L�=��IW�A�{U�ϔ�16�5��m���5����%t=7�
���}_�pDTE3�P�P�t��m���'�3��@~n؉�c�6e�����'��/��ы�]��.73�������>Sm�Dq&Y��S����{����W������iR�z>�+�Ǘb@����26�H��Ps�G�~I��K.��0z��O'nl��9�u��t/���2?=m�ȁW[WgPH��ֳ�w� ���Dj~>���m|�Z�8�	u<�Rg��A���m~����Xx���5�&��Z+ܩ-V*�iŅ�|��=�GLi�2�Z
���jJm
�e���zDl����*`�n��5�8�)5��T!hɪ���T������X�fC�c�������EK��IR�w#�F���b:l����?}�o7��N,�:��+$[��,����E`ҌYr��qP�k>��
GV�<N���� !�y�J���h����B����E�a�����ۗi�����5#L���h$��2��CM)L��T6jRꖱ�+euW��FmS���K�AI}PԨ(_�l>��g�E�}\���`{��5����)��c4
���.�y�aG��> �xSVf�C`�)�x ��G�Փ��8}�da��bk�VLh���6czc|���\�[>A0��SRx�w&�	����wzuy0G��sp�����/���?a�M��ɃZ��tӠ���:⋥f�����pde��)���l�A=�A[�bjy	��gy%��ؒ�0����8��ɤ��)Y�j^;\�_3J��,�u�&�/�j��#_�7��������Q����l+������#���ܣuN��˦��O%�t��=�[�诨�$ȃZ̸Nw;�ݿzl �.G��gQ���,�$��.������y�/��ݙ郁��`��$O��9����Lղ��P�j8�� ���L�w
�W��yN�_~,��~߸ו�����g�����j?~}��P�lA ��ͥ׃������'>x�}4�1�ZWC����!覞��in��Z�(8Dj���T�/$�����T'�R46�����*�,n$���/��z�@Z��"KE��X�l��<�Q�^����O�	�kr�Ѿ�TtG{[9�j�d��(w`snw8���Q���@jt>��$�F�~i*v�<w�mO�@ĺ(��ICd��h�*���L���G��K5F,�×�t�׶H����o��N��
U���.��UK�����b����<�b1�k�����JǼ($L*�_��{�n@]�"�^�1z\#���L�zy���0�^4�k�*�-�P8���W�SV���Dt5Z6�:~��!�q�I�*���>�:?0o�s�:�O������yFA5�ޗpS!�R+%B����l���N2�J���U�!����.K&�*R���- j�x1��sҮO��e��9�5�P�������Q�%�`a�������XXC�1��|�2y�d͂�ŧ-���'?z(Y̓s�9��8~��	�H�:�,�q\�� 3�3}.'SeۊZU�;�v-��r�7�u(_�{�v	�9]�Л��V�z^N�.&3����^�: �v0E>�N�4�Ib���h?l����<�z�L��(uw,��[=�R����aI���k�@��x[F��N�j��$Lq5�%D���|Kt����_��.R?2Ro^Y�ِ�l�Cz�úӀ������C�ӂ�>R���!���R�b]S7�m]�'�3;�����ߦAڼ��?CY�.G�3FI�E.N��3]7����e]��l��~�n፪�����ab)��Z�T2H̫��p#(�ozi�O+���^^\e c�ad�N���˗�ܡ�4c����+�Z(�� ǭ�8d�d��W?�	���L��|M���_kqF�̊�� AXS���`cc��jI6�vrf�*�_�)6؟�+0l�q�}��v�Bd��x���NY�j�]���D8�zT�4���U�:�ѯd�sԎ�C��=R���ZX�[�յ��"�un+�w3������ ��Z�7�@���X��i%=n
���_�w�=#Y�	�S����$�A	�šfK7H�9���- 憗L0�D�W�F��t�3忚A[�E;�>�R�o�p������pj^�������~Sm�s5Ɔn�U
�Y�D���.0R>�e�tk�|n{�K�S��9��(o�2�ܤG�ԅ�Ut��$�{��;��<R����,I/��/8�N.��[~7��8RW�'Z��o ]�n4���}M���p�\���� �@0��K�nu��?�(Ppf{�6q9W)��:���WzJN��5Ceф�~�;�v*1m�9kR�A�IMv��:� Vt,�
�3��oȹ�N+X�*�h���۝��X3�H:����V�����MrXXH�V�9[���@���n8I�q�sU��|�,Iq�Gk��ۣ
7��0�����~t�=w[B�zf{��u���I�c t�����L�N�2�*y#�ɲ1��o(5e�(w��>�W_i��_yk�r�H���m���J��\�����MY��wM���h�g�Md_�.��g�/�h<��9, e���)C`6as�k)��T���a�&��~޹f�lo�� E�����m�=����Qq����bZ�.�e��K'�b����5�.��. $b���T��xn�廡�#5/�YJ�1krN�X͡O��5�_G9g������UF9.^��5����y~;+sܲ=�ԕ��v��4�m����T�[ˀ���ʕ߫n��ߗvh=�̖�X�2ꄬ�[jPE�c�!�]#h�W���ydr��d<��{���^��\�=�s�{� Q��7g�V:w�h�U^4�;g���9<*�D#×	��KO��]�&+E�*4���T�z�:B#�Og�v�xVbR��r�ڭ�O$����!��C�d�d���b!^�׸�Nf.��EB �b!�9��۽����GZ;�hF��b�k�ރV����/T�[fgm�w�]t*�Ơ	�E/�KrSG��t-oIÚ�Ʋ
�Q<4n�Ñ�gk�	�?�n���̞��ʚGTO�e���u���MaZͿ6�����r�'���켿�:n��a)���%�{��0.v��3C1�pS���[���PJ�e�[�T�����ͱml�4X�Up��c�%�4��Ȏ�u�|ws.��G?���z����
�6� ��5�-��n"���7ί�>.�1b����������o,i����syHh����:��-4]9��=�%	���F8gK�yx����W�N�(]U�1���h��$甞���m<��>n�"��	,��/���pާP���I���7�S�R���g���������=������_/����\Z����r�׃�P�>l�Df�>�K��P>��}�l�����P��P���g��]����YĠ���@�U_�IYM��N����JX\�R�NaX��ڝ֛����|�uw�m~ޫHفΨ��+a�L���(������!����~�'W6���K͖����i����Z��	KM4�
7�G�D�ew�26cT��\6�K?>_6�&�=8w3zh��\�{�w`dD0؆૮-���6��Jx\���SM��TH�׬�t(mp��pK��I���I<�觺��}Z&����x2]�2A���h���'�t�����2U��ƑP�Cb�q������%���Qz�s�$f���$-�]$���l��D�f@��ćotS�:G{ۺz1v���"x�o�GhMU��in{��Pj�Zix���v!56������f��;b�6G<:�ם����{B��C�.�Me�U�i�������7o厁&_;)!ƈ�p7���]Q8�A�`�<DIz���tu~�bzZ�0�Q� ��
Gׁ�4������봥�bs�����s�]Ł?�F��ݝ.,ؾ
�،q�k�PG���۪_�����{�̝Vl�{�)0Y��'+w<��]
�+��E_.�4r�\�v�MJ��xS�4c���ކ�k-HM���ߛ�>�ě�~�0�7���"��>@[[OF�D!��r�[�1�{��b�P,HF��s~vA\�ip��)��	ye��xv���{��⫑�3��TF,w�f�*m+�����"�/�Pנ^N�m��:�p���ܫ����o�ح����ha�t�����6�H��<����s�x���C��EV_+f �C*��o�o,/�	�7�� 0%��ɾ���~�1���c�@��]���wK-ƳM��_�/S��N��Wn��G�5��@t	/�=ͭ�����U��u:T���p�+b�S��7E��7��L�R�Hn���{�0�I�.�vL�1�p���b���fܾ��~@P4Q�0U��ޥ��N^>O��#�%����+_Y�����5tL�S����z�q� ��ֹ���jcd��O�������!��-l��Q��^ �n�ٗo��aJ��)F�C�+��Ge�1 �t]�O�y�0+'w��/1n�:�K��u7��3���ͭb,|-���[��?ٮ4���|&ﵘh��Hc�1����IF8�������#�� >�����<v@��̸Pt}[-�����Ͳ�AAX��ld#yS[K#��>�V��ުXV�;�J�e���n�
�r�qʨv�;����d5���}���aw74�}��Q��\vGFǊ!�; ]��!�+����"�[��}� �*��f�x���Z�5l���F"�� $�K��Ձ!,r�,X��S��Jl��f&2a�3�xiA�c�~׼�r� ��M#������\���܎����I$�����2�C�O,������^;������dFY>��q\��*]��(��gq�i�E��x�LM�J�=�l���s����px&j?|wԂ���##�`����7g��p@�9��$�K�/�`�^k��>un��~���<Q$Xl��OV��V<���P��7��խk���?Pv�`�M��|Ym��$���n-wIQϝ02/����`A����c����Ư�%aR�&t���l��-R�Kls�������5���p?��hC坢�]��k[_�Fs<5���w�Em�+/�e	{A��[˲�V�w�>^�͂e!�y�vyw�U����4�������o�����^�CElP�@ym���i���3�wy��:����n�>Ƞ��	 �
6Xhd��q�B:�����X�u)�YԾR���(�_y�[��G�דW��-#���̒4�4��-�i��m7�e`��Jh���%B}x�T/�}ꍚ�ki�W�ӕz󛝢�k�}��!�z���ƙ��̪��ï_:�-TO[az����m��۪�D�	�O����>k.BE�l'�;�9g��4�V��b�sf��!���7��l B��T����ӷ������"�k8K.�(�|���X��w*۟# v���E��:Y���}^�Za�_h��k9��ТQ$�3F�X_r�:��︂6YEV+9
��"��*��b�����M��|�	�%��&�q{�~ݧ����<�O�s,/��x$5�\�ޕ�w�q�}��	^���-��{m�I�w�>}��
c��� 7_]!�����-|��)��7{-�Q���������Z(z��LWQ��`�?~�d�,�2���qy��h��W��q�<8<�VX}��Ï��#�u�4��x&
�=5��d�	DN�!O�ƟDs�p���j�?��;���b��޼I�����%���C��.?��R ��u�k�Ś����$�1�:��=��d^�O�{�f�G���'�Mg��I��Aݻ5O�ߛ-��4���L�A��,׋�8� f��X�ަ!Qˋ7�z���l�Hm;����'�#M�¿Z|�C�eW��V������5��g��A��?�&�g�M�����n �}��z��(q�b �YRZ��<�I��B]�w���b��K�O	U���kJen����Ԍ��K�דhd�Y{�*�?h�O�-_���>�d7g2_F��˶E����[eG�]@�
X<��/�9KJ��J�T��ޏ��/)o����
T��u�����cM*^,�"	�����T���GH����`a?f!�6^m�ƂrJ��Q���!�m^w�3~W�[��V��0��Q�;��ث��4���r?;�&���������!3���Q\�v���	j��i���s{9��ɉ&���%�{!��0�Z�ˌ���,@���2��t򷞳���a�h��t��4���Tb�	������g�����搢�?m>4�8p��}GuNv\c*H!W�I�敕D�L��>l����J���7����q��������t�n��ؖ/�)1�E��{_��0p�)P���ݘ���9�Ve&O1��>P��`�>���찬��ỹ+}u^^S���^�T���'���oo[�τ�
������ݬ�=�x���[�o���@3fO^T��,y�hn)Ё����uP��DL���������JUx&���U0����2��b�w�t�%��|�Ks����PB��`���߂�v�ek'q ���a�j񕊒C~=л2�ϋ���u��'�JbO�jFn��x8�ES�x�*��<q����=�wH�Y��5[Fr�ƨY2�����q��թ����æD�G��@��y���a~�4*��>� �>H��}���z������GL�WS��ҁ���"X�����R���3�M�i�.��\����G�?ZI�S� ���i8�׸�h���{Q\�sݢ���8�ʇ�2���]�����oE�%��I�rp�*��g�蛅�봎17b�U��S���.��k.¶b��{s�*w�R�����ֺ4�	[9g���y��:�V3f�B�Q�*���R�������ߙ�ߡ���cK�'�����i��U�/N�|l�l��f���e4���:����k��Y/ m�&wQ��=�Ш����0�ɧ{�׫�CJ>�䣣�?��G��=T�r�����Jע��H��<x��Z�2����M��"oZ�}sc�+�Jx�7ФeX���/�F����"�P�~7KKun~S���}6v�.v�C�,/��i4҇��&X���|�|5���0����V&��vr�}�ИWZl��O�;�{lN��?v�khr��S���g~,U�2��0D2�2��p;h��D�D�!��r#7h`0���f�׃ʳP��+}��l��f�E\��SS��`��_��&B	�E�et���d�Z7���|K^.Z�c$�K�(�ј k�t�;��<E�s��i���9�W��,�RT�)1Y}7�Z<N]�%l�ت��gP���Ā���춋��ţ���g�̛����;G�Ed���_r��(�a'�/�>��G�'�ݎ  �!= /��;U�%���x�m�b]�S�	nݒ��}�b�z�;2;3���z�r����-2�g�Č`n�	h������P���,�����^XN��Nh��	˛�<�c�G�|a��|ݏ����w�@��*o��0IK�J�h����ȓ���Pvar5)��}_���Lo����U��`�J���֍��7����*�,/G}�Wi��߻��f��K���hm���G��u4���SL�Nзi:�ܬ�Z{�n�����3˃� �̠z�;�g�=�0_ˇ���CkО9 d2�抆�j�n,x�``�И\N���ډ"�����'P�+�����~�����P�����|zt�C����߻ߧ|D�I��!6=�l;�!A@���o�v�T�{D��Ӻ~�gw������L���f$��vK S�b=*����w[o�:Y�A낌5�=\F;FL�N�eወS��Q���u]m&���ʳ99[��z�?]m�9���k:@��f+�	Ӥ�k&�W2�ɎxK�<��p�'��s�u���ݱ��mt�XQU���Tpl�ݗH����"jb�V��-R֎����Sy*�.F"�<O2� ���S�!f��7�%��7������?�����6�n�0�
�چ���S�mI|(S�I�����<@'�A puu�70�}0
E3��{������9�2�5	��%�&�#��0Q�(�-d*��{�c����PhW1��h��E�rP�
��������Uy�D�up} �xį���!��`�]���Dat���z1�=���,��
Y������Y��H⟢�A�t4=?���!�7�ʱ�E���&v�+u���p[6aŧ��������L��*j�f�qK=ɗ�{�ds)ɺS*�W�����`Z*Cp3������{ ��X�98Q� ��������;��^�HX	�t˧��ҫ�N��fgCHU�T��K�|�ɼ��t�A^����8B��BC6q.ݣC� b5�ě��� ���U�#�mW$U��C��_M��e�o�
ֽ�����c�ű��P���9����U�O��͔d�u,�-�4]'�|��ġg5�߶�ADC��m���Y�?b�=i�F,�G���>[F�X�$n�]���a�F�TY!܄���-0�H�fd��>��p�E���'˲-.�SEbT���Y�:���cL�R��Do�9�&ՇƐa�����g�?�7�ػ����d����;_�Si�܍��4�5��8��"���
��-':g`��;�*�B�.t4AP¹7���5=����/0�`���X�����Q?[�RK��R~�d#�|�6KM�B��0�F��Bu��d�Y5uh=U���o�Y��b��5�Y���6���%�k��R�U�[s1��(l[mC8����u�B#����p��9��D�Y����v��AR� �UQ�d��:�O0���M�]sd3-ݝ9}<��7���o��	C��8�8ct\ϋl�\_���p�4��߂_>���ZW��o�M�2Ds ��Sh�ީ������鏔�k5P�X��p�%b��&'V�$C�|Ñ����qf-��kɼ�"#�C��J~tylv&����ڰ{y#k�[��O%����6�,���b�9�tI��5TȨ]��Dm㈓�o�lZU���܈���"�����W�\��9�Un��Ɨ)�a�SF�Bq��Y�[P�S�u�_y��]�w/�3���&���m�Ҋ�	�ࠍ7*�i�|Uq�y�2x$�xbc�,�S�W���K�*:���V�T�ٹ��F����D�Up���1V��8��ږć���=�IÆ�9V�B���9���|���%4��G7U����9\x���L�M�� �Dp�R3ڱh��D��EzEt�A&���/���ſ��^��Kv���g����t�J�ov�Z&��rt�w��x���������*
�$��0��:��&�k/���,�����������"0��C*7�Ep���c���3����\2��-�@�Q���������)�U�
����{�v0���:2��H�B�luM~�)�~&{�qF@��scȥ��+D.?�'�E��\[n7}�1?�k����Ə��S�q�I�hI�/�*�E$�]�V<�ЬXFS�x������X_J��̛��$�\
�*c��~��>�㠋47����8�GLG�%?�	дE;B�K4%��y��J���-��:��n���ƋT�5 ��5�@��%��c�AM��f��_��d3�|� �GJ����z%�<E�zLY���x���b_��XY��vj�V�ߕ�hs9�LL�X_��K������(��b�v��o���(���R���B)X/��1��`���LE��}2\8�Ħ�f�1�y�KVa߆�_:����:15C_y*oE�K�Iy$.���'|3Y�c}^�F���U�?+����/W��8NDGC�N�w`����S��f�9����~1ń��?��ܳ �<as$W9έ[��ά��9�;��!'�xk�X�"�V\&�R������ƔW�	�� Q����_|��p�Ń�8jA�&�)�թ�
-�Xq'i�Oq�2u63N�vm&�5�:��ˑ��Td�,>ûb���Xw\����W����1�!Ǘ���?R3^���k ?��jKݐ>�.$LY��^:�f��  �os\D�S"[@p�-`Z"gC��������g�j�@�5=$�û()��_d�4���QΟe�Df�XUZ��U�a���˼K������ �eW�W�$�0.6t��v��]�u����wN�}G)���ڃ#�N�4�C+�RR�IL��kݥ#��첊{yu�ZΥ��^�Ե��Q���u'?=�"�ehCכ��S
��yD:�6�J	�Ή�@;��9��ߜ�3�A��� ����VOL����0 �+�Az��R�F������DY �Qj��.�(�;�y֪��������(r����}����<ֈ�z0<���I,���<-�;�D.Il�\��,����xsq�߽��5mv@>�#�>����+��e��
g��U��vUb�L�s�%�b7����{�S��e���eW/�Q�PBz@;�vq����GTK�?�����c� ���Fޥ�����&� ���Y%I��V��,L9,�Y�������y��.�/m�C�����(.i�VEGT�E���.���F�8(�tB�>�d�n���5�M��)w����y���h�Ӱ&���*���C;
�W�3㋕q�p"����ZX':Ct��l�;�3X�e|�	�޷�J�������2���s���(���2�{��G��: ����	7�.���eЄ#��(���t��B�ǣ���\��vFj!�w�u:��Jc���,�bTFJH���S��;�^ه�W*�3r�����K,��/2��0~�S����ǇQ&�iYt�+�
�D�sIM��h��h.^���JfZ��"Ub�0QR�~8��5V9�����_�b����",�#����9������E�����Y�r��,�����l}\M�&�R��8��$Sگ5@��?�����#hG�p�g_T�Rn�u�˃�?�fI/�oX�����IW��jܪ���4�����'�����L6����L����n��]�� uxO���F3A���e�57L����SHN2o���Ʋ��]�\D#���y=xB}���l/#�4�UG,�}����%m���$Y�q�c�.-4��)K�]I&W���ơK��%b�o���)���-��0-��}w����'F��M-���_�Nn�2oQ&uZٚ��,�˂m�nT��fN��W������ G�O�ؤB,��dh�UR�~]T>��
R��l[&���8J�L�3|Ӏ�x�;��Y�K�����T��>$����w3��^���r�����C�o�H:cBp�uZMR�m�>�ĭ���^��Cq& n��y��@���$�ނIj��΄����C���m�
�gM2p�<bA"��\A@,����N{�8�����e�p����ws�#�g�uL��=��YBLSkh�3����p�g±���W��������>�ud��(W������N8 ��9�pݴ��;���Q0fK	J�up.�����"��E�l/�*T����5�zˠI�TK��h[�~�H3jr����Ӭ�޽��!$�T��Xy����2��+C+�}1�k��X6�;׼�E��;�DG 6b�ɰq�WhF��w��	>��7t����=E]�I�_���8�O��"���j�b�u��}����u����A��\y%�p�+��HA��8h�/��y~��J�b�q�,�`C|��;�WvE�nI�#Sگ�-��d,��J�EBf�A6d�GTYz"̖"a�T]��g��w�ea} v+($C��J�1ި4��<�;D%o�]���E=�ƖGg� #���5�1��Jxp롷Ǎ����l1ǈ
��0����C��"f�4z�aq��ԛBf��� N̒+K9����>��rRrQy��R�g��EM&3�Фw�:J_��Q��(�Z�WB�I�@��DK_7;����?y0�m8���C��κP�Xv� M�|͕�l�7w	r��6�M��N�B/���U�\�ʎH�a�_��\�9�]���S�H�,_��z�LT�z~���������¿�7z"�]�b�O�~�ۧw�>���V{�: ��I����`Z6h���{����%߫�W&D�X6��cT:��M��a��Uƨ?�K��N`�ȯ҉��U!�����Jdo�@���)s�f�2�՞Q������a��#4m�a�(4�A�K%a��Q7S2�-2��V����9/-RNC����nrC���4q�($絬K��=�+$#z@�1y+wg��UKh�m��{�HA���S��\������{R��=@���-?Y���W���t����4wqwdWy����#5��/1�c�<�7��\��I����v�8/ƕ����8mfs�^��}

�L&�>�D6͉���,K����	LV3�"�[�/��o�'�WDG�������;a�i-*� ��lV6�t�w�lj����=�P�׫�+a�bΗY�1	߆1Y�i�����7�ԅ��obxjβX���$�����^��iE�oP����߾!W�l;X\G���<����S��L���3 �/��j���͕g�ki&�Q�&11����ݤ�F��,��=�����R�T�]_��>Qe�;����w�	s�N橁����l[�c������csYVS�|cZ�]�I,�`��]�ŗ�2�Ֆ�٩=����tTj�jS�����}��ڒbl5�QT�I��*���P��;�b�xw}#���~��_zW��x�T؀b����`Q�5,�V�0+��w�@�7�"#v@����g�<��m�qk������H��*/%��X-�\�䃢剶G伬D����%�ݾ[0��/qL_�0٫���2"�|	���H�䅲ĉ�(�e�R�N\&��fpM3��,:陖�P����ѲU�C�M=j{a�mcN���?Zث��=��������c�"�gKt�M��u��n`�1�qQ�@�p�45���_��U{oh��g3�wOΙ_j'r�}3l�r�k���п�V�0�z��;l�:������!���i

�#,�&}�R���q���J�a�������t4l<��lA>��d�k �Nu���/�:�͆&O[��X6�F̜��*I@���E�бJ\	YIH���ᴩ
���P���y
QQ��
�)yt����v�)}(%��-�5�I�t��]�.�v]��k�!w+1bX�"�v"nЦ5]��I�k�^!i�O�I��a���5��r���v��]Lf�_��om�T���mqk��JW(!��32+~�����z�18n�=�B_��ԗj?�)A��8Ѣ��}C��ZyN����(�))��v����g���cI�䶙h�u�yZ|�nim�o�ϲ�B=/'�ʴt'Q9��5/iH�?t����5�wH���y�iC�ȧZ��?�no�$'mG��*�������Q�#�h��܃�/D�aO��6|���a����5����y7�6z�P=�����[���tQl�B~Яw|�;�{HV��\�qwO��]9L�X�����i�t���X���3���8�$fVQYyf)��F.�#Ə.��1�%�O
�I8S���h�#�iN/���w%����{��D#�EЄi����}��.0ǸW�l�&��J2g���LSL��)���V�љK?�m��e�~q�fl��\ژc k�-ך�F��KA��:�����!�rfӼB��M�'�г�c�w�-a'˛PΔ�$?��ɣX��A*��K���G3���ft<��,�O�� ��E�j���0�ϴ�/B��c�m�6|/��T�P�VT;�Ǚ��;��T�՞Y�����a���>�<�\�����Jxܸ+�]M�b˻Ro��>�I�F'����y�i�ٖ��ݻ/ڝ��uq=�(��[r�%YG�i�e��fݔul�>ĕQ��j�Q��n:��>�/�ơ�;!h�Vy���4�h��C��Z��趝�df����M�=Gx�����b^�7=�/m,P��7��x4N�-�A���Q�ȑ@'[���^�Cb��>.ug����w��}����2�msYˮ�e-۶�p��ZƲOZ>�e�v-k�������}]�}=t��yf�����W�J�Z����Ș8��J�ڜt؍v������k�"jҬ J�1D4��'H�|O�<��V���ј��ɯ-f-4�|]yr-�.�n�NF�^����џ��1�t"JI"��ry��&�fQ�BDR���c�ې�@H�Y�g�_��Y����=�Qz��>��r �5י-N�;=#���Ab�l�Ma�'u�+sͦ�9uo$�/�=+��<�-nf�=�E��qVu�S��7w��P��2����bŀ߻$�����_�\碑�0z�7�(K��9�K"���Z@Jz�$��7`�f
,?9gLq[ �1�=?F-i<�N
�0����*D�!K�P����K S��x�(��-�x� l	z����B:��6�hGp�I���\�6�*�t�ŋWؼp�0����p����V#[�����~����w�#���V.M�i�+n��'g�T?v���!H ����-��~��e��n��Z?m{}9�[�X�J
P��"cc�&7��+���U�3*���=�Yi�a�bQ���HːK��i�e_o���ab[�+����H�j�hX�
Zת|7��9�����'N;Fb�.�ї�١:�|�?o��R,\;��#l��/|=��e\ڀ6Ji����Bv�1�1��x�J�����X
��!��W���ڗW�0mG�i���d��Qn�J1��Oo/}�[3���c~�� g��v�l��T������677��ӕV[d:�w��Q,'9��#+FFJ��Ł��v���)��4������֘ؓn@gJ������n�fD�@�ąO-R��w�F�f�)t�~^,&�9{�gi���*�z{�$��	�Y9�`�^.����6)�Γ����/��6�bY���*2�<�M)����A��9��_�,��
�[���*j�HC�8�
�e��ʪє���&8u����w�nnǬ�2=��Q�젘���! ��������4qe���
��JS%Ry���٠�n�	M�E-N^E*��&��9YH� KO�\�5[�dFo��]w;�>W@�`�*�F,� �[/_Z��U���&�b�}P8q����|黂M�t�uK�0�-Z��|��Dg�� P~���pC0��e!j���R"СOW�q9n���,XG����%9����%y�!O�`ȧ.=Y�uߥFB�T���͢][���~��
���v%P��c��F���)zs!�J3b;��/:�����^���|6�i�Q�] Vu^C��v����w�^���v.���\��j-�i"��9�8(��kn� =�p�zE���!yo�7�=3�'z��dm1�I�9Zm맅�����!���%b �5��سf�=�*N�n�B�p�(��з��h����9��goP��&���*I}n������r`��~��r�!��?��¬�G�r��Q,��xɣ���U����FOm�Sȷ˳���N%փ�b���;�����&B��7S��=]DL1#
c,1
�6Ϥ$qc	�/�7�씾������������ڲLkf��������ʈl�'�u�UK;ᤦV�1�3���� |q�!���>§Ί�����j�j��}.�v�g�P%��b��$��nȗA��gE[򋺋�>,�9f���T�����Z��1���?�~+�=���|CL�������'�3�cATIcq��\�vDR�m$������p�KI�!~S-�"��r�G4ם����jiL�^��<ۼA񹸑Y��d�%���C��.g�W�2>����ǢP���lቌE_�g��*>�?�QWJ�"����u�-��|FY�p�I�΄��(����_���]�N�U�<�Hh8�HJ��{�餟�1^�p�:�L1�)���~O�ǁ����h@�:r��|骃~�� �Q\� �� 閽�si�Z./bP&#�">b��U��e�o"�JIΈ�SE�	��+�=&"����eOF�sQ垈�S�:y�9;�ritc:4;{���L���&������[�q\����z��(�;���V|�գG�L������1�sa!	�YAdl�ƍ7�+�䭡����SKm��� ^���T*!˂�����ѓ�r��#���f�&>EذE9�%M�ɕX�<��Y���Gܾ���K�B��+�tH����e�p���:\�
[L ��Q����Z���Nr�h*!&��2��!�u�H�O��ݎ�=���1ߧĞ��P��+��K�	y�3�U6��r���@���������eI�]U�8iւ~������O���[Xw潇`����j���zS���w�h`�aA�X# !;�o�tW�����o��|�J5�J�X��ţ�V�� ��͍�;��\��������@�e�c`>�t���,�:h"��kOQ&�sb��Bv��<\[����|�s����b2xH�O��� $_�!��f�z&�9�%�CՑ�=����*�U�D�X�y�̶I��D��ܲ��<(C�m�ru{����&�z��Y�Z n�M"��-?�F}0�	*���;��m��jk�e�2zu��m���1�'��dLF�$�k��iw�>v���>(����le�(�����N�W�I:�a��}�Zw_����ǳߨ���zզ	Ī��D���&�������i�*���SdL���\6]X3�Y0���:n\�7��Ϩ������=��bׅ�TC��:ji��P�H���lb���� *Ɵ���)уb?&�(E���|x��^�OG���LZYHsl�VBD�P2��|V���[��ǒr�G�M�R8M�$���\�P
�����v�K�}K�-�Hn�NFcGϚ�J�V���37���~��O��N�;�����.5$�+��c!C�BrT&�97��\��iw?DJ�ݨ��>)A��U��+I:E�i��;FH4�&��E��0E��;��[D9�`���T�5�oD��YT�Gq�jM����,�F-%�7bj�+�%ʼ=�ۤ~ޙ���j�_�Y�_�\�	���;��t�P���mἂ0��T��#�\�����GZ�H/��S��!���'�R���1�⻳��������pX��Yk�R�㟗���P�%Ԑ9eM�l���
,� }��N��/���$t]
Bwi��H�~���Ty˼���[���v�B�C��{W���T���X�
[�7f�B�7���3T�d���l M�&�%�gs�UR_8o�Gz}V��]־��$o()��O"��j�-,���yƵR?V�CA�95NgW����D�eک��{_Ʋ��3���#�����kp���ӣ�������+#:5ӓ5ߡ�K�\�T�z���券��X�ɉ����h,����e@��|٧���\�)����2�^Ey��"[�tP�Ӕ�Yt��.T���HT�t_y�U�A�H+��zN�%�^Wy�h��k���],+��N��@GIt��,��m��Q2���cz���i���[��U��ӏ��?�~;�NZ�|q�r���q��	8]# �J�Q��cY��g�������X)'�;���
���Z����b�$��w�hL�)"]k�6������i	D�\I�L:�����1�Tq[� �m��Qc��Z�t!�^�+7��(j3�aU� �ijBK�ŝ���s����1И��C�}��L )+.e�����=,���ji��������\���H�X��r
]8-�u����$�۝��d��,�F<HS����/ͭ�t<��f"��v�^ V-w)�~y$'0WFp��~����0���}k#�ۃ�>��f;��r+��z�i� `�O�|'�(��ff�	�(Ѝ�yjBT^�#: v8Bb�b�;����ʡ���z�)T��Q�?e�H�.��=�$�$u�44|4"zw��!A�.�UeQnRkml]b�`��|M�/��}�
YP�X�#�����c	7-��a��bc}To�����ē��.��� �JUf���s�K���^���X'}�%���w�Ͼ6/�Cs%Q�/ڱ�e�eH��1E(N�m��>��������e��|m�w������xo�o��8/�-띰���4��ÿvo �?�d���VJ�6���t���x.5H�"�@`	�?o�1%���.;5{@�.�L�C�<]E�>'���I8�ޛ� ��%N�P�.M75���[�-|(� �Fؖ�J
,���P���Y�݆���a�f
Q�-��q�����QC���x�1�Z��x9y���~� �Y��F)Em�y��f�QS�ѥO��Ǣ6�7J���u��&f˺��§�;(��g��a+��M�fYwx|���mT�)܅�@F\�B�W�O߈�;�>Z�J���;�a/��R盝�D�T��������Ƒ5޷���'�R��=WA;C��<� R��j�Q�������8#�1�
J�^���!X���n�gtʳ��|NK��mS{�[j>�Jў��`��9�Nn�з��ל����^��X�oԣf�"ڡ0T���� ����A�I1�X_nY��օ�����JX?��dQȕEq(�j���;�d֡�#5�#��*]�&�Ί��iӔ���Tr/�&;�5��L�2=a@�T|Dd5��d��ݼ�����D�%	q���؈~`U��^n)I;�����g��6�R��w��p�3�¨�;��h��7�̈p
���]H�lN/�syy���U����[Ma�@�7R�*�ewZ��yd�~	����������1��X�y��GQr����Z4ָE,�҂����H�p.S���%��@y��ᑨG@5{�d��V��ƴ)R�?M�94��r��u<[��L.�N9!@i���D�#�8n8� �n�T����D�Q�z���??[��R���[~蕩��V#�d�4�6�l����</{Z��"�2Z:N�blB�$l�O�欖�!�MQ�;�u�>$ ��ǳL<��d��'��?=wK����]�[9#��b�a�����p���C�al����\��A�!s�uqD�n���s���͓
��S���n���@�P�#RT�*��dw�3�?�ǈ�p��ׂ���_/�C�-q� �~���'�b�'��C��W��v��n����7'K8\Oi�a@$"�����BaS@V�!������+���s�	`��e���j�|�&o-��5����Ú�Z����^!�G����V��ĸ�����8�{P+{z�K����s���Ŏj���f�G��-��?b�}�Do �Q�v��Q�n��|є1�q� ՛�����X�`�;�ލ����[AKC�(�j���5��K�Bj�~x�j�"}NF[�'KM���<���3��;�.��b�����p�2�ְKP���K�Z'��bI�m7fme�UH�Ylk�4	�S�$#:��m�d�;�aDg�^�SU��fJ�"X��˴ 4���ۛ�D(;��o���#[u�c�(+��K���V?ʈ{!��W#�z���q�)�]�ҥ�(���kt�m�׏ ���M?u�oP<�'��g�
eWg?]�_+1�a?���D�R�Xw���0��	[��2�����q8���_X��2A
�}��%������0ۃZ��U=-�����t��j���v��7�l��K(��reOE���z*�Ez~��E�$����
����c�d�6Y����(�W��q�o��oƿw��y+�o/�pS�X�l�u���(�T*��[�{KW�$��?��8���6�Գpp�T;"YۗJ"�xc�N8Ҳ���L��(��k����_p�cjس�E'�������`���.���ş��TfQ�Z��7�IT�e�k�R���nF	�!��ླ��;�bg6 !��6�>�52��AVa"cMQ�Ѯ�`�D ��I$��9��3�!��Ԕ'�|�=�a�����S��G?��e,M�C�kv���rfA�,]��q�c+Ŋ�+�*h�c�]�#C*<`"�����="DO�?>0��F;QM��2�lP��X�#U�]�W�h�=�Q?���^uf��	-��VGt�r]������򹃨,db�>�J!$G�����e��<��HyS�Όh��Փ��T������i�[͗����?.�����{�Y-��(� p������+Ǘn����L�7y�1t�-y�2 ?"���"��M�
�&e5ŝbqe�5�	�ҩsl<HO�Fq)D���cf������<��#Y�
8�dx�ŝaA��oX�]�e����h�J��zᬒ��.?n�-5{���$�^mݖ30�6)ߛpa����ʀ�L���k�U� J��9#{�I�%�H<�9"��R��=��g�d��S� 7�O(\d�h��D��[�#Y6z3��H��^
��;�vuq4{ߝ2&�RZ�m�"8���i��j���i$5�l.Gq;���0IY�����H�=��H���?^�L�t�r[9��V�AA�I���s�J�i<�P�ԧ��?Bl����^|� j6�F��t_�E��P��|f[�M�H�����wD�-�8�c���i�;n�@�܏-��b���bd^MM��Ld\�1OX5�B��%6�a~^7�H�,z�CN.���dB�.�^�]zVL�w���r���=��vNռ̚�	�t=���B;�X�Ք��! �c��y�S�f��MG`kx�cz�H���L�D��fȵä
%wq�ϵ �˳����mH_s� ���� �9kh9ZQ�"wC�/q �1��/c˜�!�V�����O�ߘ&Wh���u����>bQ�Q�q�]�����dl�#)�AM��v���D�[��Rډ��Z���#ԣ�lc�nw�_��t~�s}[,���x�_����đ�ѻ^�Uő+D��6�'��1���}N痔}�{�܄�;���!^}���cKMv�Έ�)�����L����=L������:Yb��ZT�A�9B������q����	]7���=&T�ޑ>����>�ؔ�[�^�il �K�#�٬�%NF��fA=���[��`����@���{N�n�V�Q�ݶ5㢯�q�\*� �/L0Z	R�F�zoV9��n��ok�M�Z��w�Z"k���F
�N"�����m�<����N\�tr>���=��[�Br.�
��=��L�g$���b��ى��L��a�3�%n��6]�vqA�� S�&Qx��jD
�һeA|�,�;�R�:�j����zJuU�Ka#�	��J�*Upt9'esȸE�}a�Q���t��{[���<��� 1%���A�185�Ǣq���|�o齖g�7��/+�x�-��j磈��'5&�c\��ɗ����E�&I���M�P\�,�M[�����|�cݓ��[뫮� D��T̢h���y}lc�+́�#?��I6�GvW�������&'/�tv=9�K��ueڨ���"�����O��UT����j�$�V�������A�H��u|���� �h��<(:^JO�(��= ���x�M=+�ɿ+j�<;\�P>���e���A�[����:),��fiQ�J������-a
q���#%o	�>쿖75
��0dȍ�$�>HMs���<!4~_L��	���]�ļ�I��p�KS�(�mSp����BM�s�0�����k�/
-xofr��,� S?����G���7g�w�*�i+�����1�`=bJ�۾ۨ�ǧuՐu��+�.��C���z���ZUYkX��,��5����o��Aw�-�i��!�����D�WW�0;�{��Z�W�Rk��.�8�	-��N 	��~&���e!1�Γ�kz5@6C���R�]w�o/krl�q�pB!�W��y�p�oc��1��C�n���n�"�Z���HE�b_����i�!#��f�G!�r��7[���ʀ��ܢ�Gi�o��`2���k�91� ^eok���ܸ�Cb�	}R��~;8t��ø�k�N����œ}����J;#+�>�����.��߻��q����A���2��K�^/\��*%�t9[ٗ ܚ�_���J��=��h�?IOdT�bG���
en�M�	j����\�0vN{�>S�>���~�h�l�O��	X`���s���5^WW�ajs��=���{���o��� �!��Q�ɷ��Y&���Y�BM%O��8��<�3��+[n�`F�+�RF�ȭ�����$�������P��&N�}R�����a��J��]�|s�K�a-�}���T��-ff�!��������;�*2�ߓ�Lo�l��{�F\�0���-���36�N�R&��h?$'�mj�
����X�*�0,��HT��ؕu+N��B&���|�M�s,�}�.5i��cfxD��4_A{���&L����dg�ٓl9{1�{�?�w�(�e���К3�����(<F?�E��B��;Ɲj���-QP�}���8�	B�[�J�?�,���+�3���T�5�E�"8G�B��$PDq,>�=j��w�	�F}9�����'3WȏL�w�!�M���8���y����������z^kN9,�]�[�0hTB4����[������8�:xY�yt���Y'���y�8�ϹU&�4�6��GD��D1�խX�}��BPg;�[znҕ��8�;#������%}��L$���&ڧ"��V�Qi����9t/�T���%#=�Pp{��j��M�x�]9�j�႑����z��̩�M�Rmr� k5G��o4�+#G�fԫ]�X�p.,;4��`�`;�V)lq>#"��@D/� �ܺͧd�c�Z�g`/1F�d��۟��=I}�:L���r-��	��pF��������JH���iƴ鯃�:����72�_��tʯ�c.��*;���T%za�lF��8��j�f����ʽ������[q���h ����S�M�
V{�7*B'Oj/�A�ڙy	Kvc���:B��)	�t����5k��f5oi�r��ߐ�2��\5�Z��UŵO�d�~��\�HY1[���v��4ХrV-H�eB�A�Z��p�,�s5��h[�ї$s�reU.�)����W/��];��YŻ����������m�8��,;M�G�h��2��j�\um\Ȅ�AW"A�^0O;5��^a�"!Pԩ'���-'�OF�
&Ѻ���si�I�$+�z8#|�LB��rٛGϚ�p��G���K�<��3/��l�R�~�/�v��˚�5r2&�ķ}Z`�c�mr�$���;�8FXC<���B�� ���48	�1���pn�\4�@'I'�:�xm���
�I��5�����fE���Pn��VĪ�+Js���NRY2l�{��Q8��1�������(������9+tE��e��t��������g��2��,��_�$¤��".wA1�c1�3����3	S����M<ӭM��ܖ9�E��	�y���j�FP.���׻�Yf�n�y�b�@���,S���&������)'�vW^^���F�Qi�?����� Cf��'�w��%_���w	2�<��*�c	)�qU��mLL�}����N�w:��.�� ��<l���
�q�~��
�0��KY�5c�}o��掆��	;�ߐ��_���U ����X.���pro�vb���*"��f�-�`*��\�"U���I��,H�J���t<b�[#&cSu�>'��8��馐�H�hyqK�4ب�C�r��V����F�֍k�.3��1�\�[l���cL�<����dM~,�;��^&�x�q�Q���_�����	����_x�0�������.�DE��-N��e��
����4&c0�B:W�sm&�c?�	��+9*�C���]I�����y�@ktqW���"�#x��4�Ƞ��Z3]
�{�	���ht7�����:._�jpis0�J|ǥ���?�PӐD1�N�؉��w"���i��v�����\yv���Uf#��K�H�Q|*�B�D#��x��[;n> I��l�c�Q�b����7v�u� o�d8�) HEE��-�S[[]XH��綡+�p
����зJym����-�v�澱I���BG��+a�۝��ݘ�ܧF�*I�u���S5�f�->��wIf��Y{Uu|��	 8��<��/��B��;�ҏ��~�>$2+�O!C�BF�)�g1rƉm[�x���G\�6���Ѿ_^��a����߬��2�$]1g��2,hU�ad�%G4�f'����&��>ߟ̰Q�R�0%Ԃd'��m�����UgpsI-���w�q�v�+���Ƀ�&�X,o���~Zˣ�h��B�Ѭ��;-��4܄~	i�t�ӇEԹ�_�9>QbNj���v��n>x�u1a��hD��"}�_�U�F�]=�o�4X(���
{�e:J���O ޯ��<0uEK	���F�ݥ�;���6�!�����L���.�M!fL�p�/S�@�q_z��E�?��J�-B�HaJe��oe�.�>z1��a�#zNT��$�@C�hlb����i�D��AmCX�MV��1H��9���Ba��<0s�e2�0E�V�$/�[���c/������A�)���V�w��$�|��6�'��Sy���0)�|�����/:#6�~�����{��|<;��>*4�H�=d�#�;i�����~��U2�4(M��d���>!������Io�4=F#�V��٘�bZ3Y=����a�ph�.e܇bu'��cmm�#U���%Z���"�p(V���Ru�.��KٝΜ)�ƅkD%��V׺M�饤�o��<=љ���o/���8�L���k�K�"�rV(��U����1��L�ٷ1��Kvp�}�K	k��3v�~��b<.ɷ�NKɮ�ɝr�� �:��y��R����=��������_�cL�7w_��=$b�<z*�ۘ�w�>`J5�*�k�y 
N�a/A|q�Fu~���4���7�)��!/��(r>b- �"�θ�M~��"�m�5��n��&�$�F�F�/��5���*K*lD�m��Ѹd��n��X�y�� +����'ȴ��%�(@��SM�ᣟ~%Ѷ�@�	�e��@���4Jr�T�����sǜ��@�R.� ��l\.O"6�[��!sy��(�f!�B��2�u��\�Ax_��=7��G`Ō�.�C���~��ˑ~�Ϝ���PZ�����g�֒SDΪp����$O��/ z���D�>*���@�M!E/7X�A03�(���P&q�5%n?��-��#�����U�$��<��U0;Wʙ�q�n %�z�3��e�B�TZc��n��4����B0Y��
��*��A�#��	K�U_ �c�e����J������a*\��&h��ţu�Ҋh�/�����m����)��_U��'����H�?Fe5�a3�&sUE�Ap�"X�H<
,ä��Ǹ�B�㔛�TL����Q��;�2M��I��f47"��w�&:$r)ߜ�Ps�]���[�=Č~�-�h�[�C!f�O[�WI��������d������R�̘�6�;f�ؾ��]����68�W3�qW��+�������D�̏��>nn�A%�ܪ�j�!E/�+����г:D����J���?���Ύ��N;������[\�%g�K�[�S		g8���#�@��&�m�w�����5�	G�R	����ͲiX���n��xF۬e9ն-뀃�!\�3�<%�!c]�I����(A7D+l� k�����g�F�bE�!��zņl�kk�TpC��d3�odY�	a-6?��>��(q����Yn^EvnU���$9c�q���y���id ��l11�6��e�ǯ ��+}��~s�Q\�'���*�fF��5c�����6��B�0<�0���ި&����MA�,7�0`:���˸t f
�	J���I'�I�_i�/u�?�X�O�_hL	�&�H�~Ԡʝ�s�V�� q�<F�(�;��S�)]P?&ΐ}��?��R}S����嚝X�b��}��
�ȂVP�vO ����@'ogaѹ����A�f`%�(nx2u=��L��R� ���vo�gЯ��ҋKA�E��Υ�C235��m	�*G���Z���W|��j��h�9$��ؒ7xH����CT��F:_���J'ibp$ns�{���Κ�\P6R#�*�XT����R�X�ܟiO_}�0P�i�X珣�\r��'1D�W����2�0t�ԑ8���i#&� ���4�%��1�U�4����-���
z5>ڔ�jJ%c�Y/gR�d˱F���������%��)�\�6�'����2i=�*��G����ȧf?������dz�X�j�İt$�Wia���1��l�|���4+�]e��
�lE"ω���ߤ�[��c�%��B�L�Gk��A4g,�f�9���O���[���,R(t�,���zHlDj��4CYVΙ|��T4>,&�<�jKa�˫J>gG��GDֈd�X���;�)�#��{�%:�F�CP���]�g �~�e�\�y&�PB��&���B�[U�1c1�ڌ2#ԃ�Z�ow�I�z�Ɯ3��,T	�w��O�-�L7��h��,R-2"�>��Ȅ9���
=�*oT�K��찒:c��k�5��SN�w��o{���;��
z<�u�k���(T+���<���]H��:��+�p�C�C����>�c��c͇E��9�y0��P�{�[�.>޸CK���X�]Vf��i�ߠ�3]H�rO�ˈ�t:�z�5衡��E��z�|�.s��w�6�p�	b�i9*���
97u076��P=��qի�c�e�I<z=Y=��'N�t��]�v���N���e����xf$jH�<�yVA�碛*O�����ǻ.^�*�7`x��$r��铧��2b�&O����Mm���Q���tV���
=u#���-é��N¹̇�D�����_yՀ*!�6�������Cz�[�������k�$Vi�+�|��f޼vO<[�ѹq��`���`��i<~5���%]�����������2�b�
d5^�.���l����ľ02;�A�������[���L$Q�+<�+�?n���6�I�d�+����$r�{j!;�~W��v��#�֒��Y �x�F�G�f�O�d#"s'�ޘ�-.��A_P@}����.��O ,��l�v��2�T��J G�Kj�����H� u��Fne�y�e�dj#����^�n���;�.쩮���/3�@�Hm�Z��p�E�?x�4-)�l�4@�$�Q2�H�WT�j�+<j�[��@%aڲ��m��b��c�Ϣ�k�s�9�z�^jE�P��R�c����1>�d�u�I�Gj���Խ��_�e�^>�%�kD<��iA�EJ^����xP:8𳲓`yc�A����1o�q���zC�Jm��� �[r��Tl~D���3�oS�[AG�_�2->(��0/o����B� �a�*QT�ϓB�R?Rr&�x	��B�d���@���.��è��G�p���V��.��r %�0*T���.W�^C�����jEݒ�Ks�+�C�m18����{���;��-H?�ڕ���߳�%/e�x����E��a$���=���k�Ҭ�V�ԄO�����}U����l�<�}Y}�'��*&�*�O��>80(v�^����@T?�L�����c !��sQ�tJ4|����jc` ͑q��K�arwmƒ��§�K]8��k�.��MC��?|%{#Z�������GVV��h�T��|������!I���w$�^o�K�:�˽�a���ɝ<i�c-��q1�ë£��9z�WB�7S�&��H����G	[y
py�8�N�c�	e�7�&N:bӖ�'N�@}G���\);:�_?yW�pr�ǤH9E�K?�Z^]�\}��͋MT�&)��U�2���x�Apۯ��?7#y���������k��7��Xf���O=L�J%�S�w�Ȕ����*��O��U@RZ�t�
M�L����*\=��d��c�t��K�v'Y]��u�PЕ��1c2jR����8Q���6��l��N��H���)�I���s���Yʵ�<9����݄c5AUq~��5{Q�(	���Ec['.�hI�S븓\���=b�-�9�F�ũz��h�
���{q˖Ė�1�hF�����k��2�Yw��vݎ�����@Wu��̹dlk�r=�=��nV$��c<��˝�Q��\�]	tF:�E���[�yS�2�?*��K)���%n�%�'N-��|�����-X����M�"���RQ(������|-��[�s� 6������j�����"�>���^��+_�T-;p�"B'=2S\�Xl�U���x�X��>b��jQ�4b���B�1���$�3C�c�ͮ2{�'e���N������2^,�?��B���y�p,�Ԁe.{TiIN_6�W��cW^��OWo���}�'���nMߞ5Cւ�|(|�{H��� �^^;�tqxA�Z�|*�D�*1x�u��L�xf!d��\�OKע9ހ���襂��\�+l��Qf�`�䃋���~��-��Xo�9�>���4�o+g�]�<F�G��U00d���i&#�����\�@��p� ��n�U=>�Q7}��K���\}�rO�<B�#4��*�/�Bsq٩�: H�R>��#Kաxc�� ��p�2�tk����F�8WU*N�M����>���eFw��������i2�=��W�F@�g)��V|zl.[�I��aL:$S[�=)��*�3�j47��|{��)�49 xtfm�S��p�K �<VC
y��O������"�*d���9�mR�$L���?tYdj�����g\�N�v���P{f�<hkF�,�[�}~>4y�o'��G	�d��������9?`K�ч]��Zr1�*�1$�p/u�� H�HK�ިǀ��H��1o��.�P}��W���y��k0�,썿M��k�ݮ��r��C<��*p%�J�;X�t���w���Y�m_m�6u������s�(Sq��,�DxY���ė˒��8+�nDym�g~
�Ꞌ������Rc�W�!�� -���h�M+I���1�������0�}v��N5��K8��3�Y�T%��6�4
`o���A�g��,�7�y�z��)�j-#sD3�-:���~a��lkfO�ڲn�.3�����O1�]����P.��]IF��/0Zۃ,N�$t�L&B�U�|8'�Q���Uv���,�a��)J�O��0��ǥ�aX�)��>놁W��z������s�W?o)pl.�)Ȃ�dU�����S�8���&zŗ����Usk��{�I=�v��yq/s˅̏v
d��O�Ϗ�#���3ڲH7�N�8y}e��:.�R�،i�C�E
S4&�i�P���A������_�trW۱c���(ZC�%e���RxtK8$jG;�X­��q�a��[�jq�J����U��s�!���'�q��W�����9m�+��[�qx��q�[���_����L�|��"兺bKx�)�lοO��&�Eq���9��:��^_���\66�$������R�s����3\�����d�Z���/'~�+�	���'c�c�|[cj/|Bh�L�f� ��o�ё�������n��D���CXGo���%�kk�*/��(��t<�5+
=�lmb �H�,�V��jp7`Do��Z׹i�qڊ����޲�O��g�s+dJ����g�B�8Y��-}������i�8_�����j�lm����%ֲ�D�<�0�!���Sۊ�C�0����$���":fD�MH
<�=(W$Z_����|N6�[��|K$����熄�L�~ܢ+�G�pe��~z�Iw�$Um���Yl����ĞQ�0gL���dij��A�A�C����q�;g�����JVSՏz��`�x$�D�8]�!:4	�,tQD��J<��P�Mr��~�5#T�ac'\�{ƜX���ߔE�"�9�śoi����>�Z��,��%�8:���>�F��h��.��N�l]pk��3I�k^�0��#i�5�+p��R�ʅ/��!��!�Bk����g����cϯ�w�MWl�i���.zkbn��J��'k�g���.]�����_�����S��7ľ�У#j�	�>������#����U.��E��vf��Tx/���s:�9�͆F#����8�ݷ����]��w�>(1H7R-F|�Y�>�	�5!c��*|�-EPI�M�f�9����EކJ�lX�iM�?�!�"=kV{-���1�lM��ڊ� HJI��(�0�D����hƐ.�!  -a�]�����h$65����y��#��|��jw5��݃sG�&�Fxa���|Y�OpppSK�z ^4����w���^��C>_.i¸�'Y���a2��M�J�3RƟ
lʢ.���Kw>��E�}@�eK�8a
���=jo�P��β������[N�.W��I<0����-�o�S�nw]?��oN��Qa�$ѵ �z�CM�c=�橝�C�?�l������x��XdBuF��dO� ���ʮ��S����2mB�1��z!{�9�<�U,f�ry�Gmn�����=pv��ҡ&�ZZ�!03r����^�}`�I$��|7�,�������adav@�����,q�b�I�Q�9��!��i0�&����3�T|���֪,�(l(�a�׷���Z6W�c2~�\v��<�uN�P�m3�P��x���.^��-�R��p������(���$�<G31���}�wX�������d�[�w��Ye\]�:;�Ǘ�&|R��R���$��<^|�eVmo\�v
@=}�CkR 7q�� 4��y<� F!���[��ǀ��Mטg�u��A���+��&;~`���B:��������{���D�3,+���/�lY�k���O>2j8���jfM>��"Ʀ���}\|7�~`����o��صJ�T�����v&���P��!�#���[��L�m�;���E�׊h�^/_L�z{�l����JW7�h�П�}A�ɬ�8QABuD�#���wj?$jgrO�88�k��]�E6��zہ�{�v�N�[A��� ,�����.�����a:��8T����[k���/��������,���|�D5t�;������5ʸ�8����O4U�hv���O���O��ws�ӛG����~��r�Tc�U�ˇ�����EM���1�W��1�p0��_]=���bB���ǆE5ޅk!��8���So�8&?Bet��-g}���B�Y�7(���k���G8'�Hz���`1�|��T�N.���"���=l��U�U�ev���튒m�U���D���&ۘN��~�y�P�0f3n��K��O�w��=H=ۡUq��L�5ʞO��|Ap|�;!lqѴ4��d���1�'H�'�f}�Bј1��ΏB���M��
T�%�}z6䞧��Z$Ľ�>D8���1���Eo|Y٥X�(����-3auC�?O&]�F�z������?��OL�A}���%��4��w����uͯ��1�)�hSM�ɧT�詤�!���H]�w���nݐ�����$y=�3b��6.�:ﰛ��	���]���,�"�"���J/[��z~#����Z+><!(e�g'�_�">�\w��fY�s=N�,;��OqkT�ED������*/-�>R�:��������'��||��n�D�%����W��%��{�1�Ӻǋ6e2����u�'�xR�#����F�OM�0)���FɺM2֌�H��2��υ=8@	{��S���,���t�ƗO��/q�c��y�(�꨿9̋��;�Ox�Ƕ[8���z��~-;�A���u��Ȇ�x���_�2���:�W���߶�]�
_�a>g���=&���!¹�a��=j%�
��Xch5�q�;�����}ZZB�A�U��W��4�ǟ��X��s("e�1��Z�g��R�fj	����xܢ�	Y�=n��{�Q<�Ř?w^�����Y�vꌝ���Xԕ"߲��>Z��X����םi^4g_%#��������X����n���t�.l����W���tW4y���8v�ˊk��&|�:6Q��8Fυ[V�|��Z��H]�o���~>�ѩ�>j�������'AWV�h��	o���Y�N�	D�������
[���2{��n�]�	կ�Rg����>`�l�,Ռ-U3���/�V���x�L.l��ڭf��
�8�V�"��M��`r��|�{|��)4�����G�g@V���Rv�d�ͩ" Rr�ѵ�'f��%%ER���tm�����f���Tφ'�Ȱ?�.���yQ��ه�V�(Wc�Ei�dD��+���j>� v*��W��x�R��3��/��zc���`�L�g4�Am�3�;Ǳ�w+#ьx.ɯtMQI��ǎ$���_ĉg�{cǸ�Tn,��_ӎͻܱ?<�������@�ٌ���4
�Bg�c��lytl�봞@�~`A3�2��ZhY�	�=v��X	�Dw.�[��{#�ʫ�����RR��%��|:�J08��8hg�y}E6��[���xU7׋�XX�Fժ�q]G�%N+��UB���lڙ{��[՛؟K���e��K�痹H����9j�zV�M(b�h�f���� ��;��-0`C���`0�p㴃䳗�c"ߩ�زG�_�2�kk[ھ)�n�O*�]��������5�͹&/�&��[��"d٦x����m� ԃ[KUC��W4���ڻ#8NL��"�|��s����`���H�OCθ��Tț�;iiK��Z����ב�ф	�Jae���ڶ��,�J��Dk�w�[�-l;�1��/Z�r�rߑ���c��ۓ#������)�yG���4p���K��U/�`ٯ�	�y��84��w�>|cgV��4f(��������f����iF��<'kN+'�a�U9&���eI�_�(|��N�I�_Ϣ��k,>*��A��)���
�A*HJ��g����9F��R���и�X�9�ܟ��!�d�Ki�V��d�CM�"�ل5��%��z�W�&�n���f��PUv3u����SKh��������}����R6����@�o"��S7��ν��=�DJ��W˜��X��:H�3�<�<���o��$��q�ozR�H���s=�?{=N�S�}�Ѽ�~cGUy]8�A�A���-zD�/P:rz�ί)��%Tи{H�������d�1����Љ�P��ԧ�=?c�����'������7��G����<,D�9����,ܛ)Qu�7��s��/�7�gl�?�dss�!�?�Y����2�)&2jKsF�{L!q�����Ј�6�����3.%�`�D��X��.h���Y_1�β�#ǌR�~��TA�	��������!�C�$�J��y����za_R�#E�b�-�c���ߚ׌�l�fӛ���Z�+?6�a�/g����Y��cETx���9F
'd�|њI��/��M�mK+�[�"����>����{�_K�UT.L��]q���O��Oծ�qa����Y�꫾W��f�}��O뙚��+B$�f<9��4��Z��r�LFO�7��9R��7�G0��ϔ�ޏ��F��_�����>��x�h}"1��$s�|��s��fׄd
=�ޙ��DWr�P��V�`TE�%�ޚS"?l�>�'�K����K���X�M���C�v|�e=��e���ʦN
,�z���#D�>+<]�Z���>"��D=>�hb�P�'�m����%���NI��>��-�ϣ�y�����9�jN#��$~���6��C�y�nT�
1�	:\���2��ޘ�s���k&&&��k c�e���i6f��߅�z��f_�M^*}�H��^�A-�G;/���p�뢓�9�ݑ�i��(W?F���-Y�� �mC���(F�qL(���}��_�I'?h�#��'��^�o�cY=���{VgB�=����v�hQ�r� 8^~�W�3ZM���q!���>r���V�^�z��{�7wk���B���uA���A=h�*������5�C#l���r:�����l�����.�X~�m ,P:$�C344���ixI1�W�&�w�:em�Aƪ<n��1J��B��%��֣�A�r{wS��",ﳓ�x�=Ds}�xn������i�#ioG��U��a�u��"�x&zھ?t~HN�(��gן�:�y�d?�ȇE��ڝB��P�O�U iI}�Wp>��j�Whk�Α�#��C��L��(v�+�������1�F����G��������l�zy�wt�f��Y�d�ɩ�s\؅қ���I�K~d:.І��/���X�NK�˕V�*ʮ*e�7�F�;n_)�6�_�����&U1M�Lx͏Π�������\w��B����p����}���� _29~�.➧�9>s�Ys"�v/b�3,e_Wع?R�o�'�hezB/�� R1i�s�|У;(�FתٌX��̽�^6Y �ޭgk6�x�����ZC�/_&���Z	�k�i-~�~c�N�v�k�R	H$���Z{��+*�G�����蝀x5v�Z�U@5�GL����K�oE�?�������&J倃IK�Y���}(d��%_���^�`&7��b�A�D�L?1�OT�]8'A�n�+nr�tS*�_��T�l���������7�FC|6Q�������U�\��pN�X��Ӂ(T6P}}a$�_x~ �i�Ғ�H��g�1����֗�k䓷�hu��R;�4_'5������:/�עo��I��L0u����r �vr��" Y���8dߪ�/�v�|=�-��*�E1U͌8j�y���~� ��/p����������~,	0�
�PY}N�t�����i��3f2�b���!�"֣4٭v�duP`-�\�?R�r �C¸�ФT3o����gs���� s?�6����X�;>4��Bv8���:��~�1�t�s�ȍ>�cI�᪩_n!��)(NمX{��S�I��JeQ�<#��~Hi�;S[G�eO�.��1L(V%��q6�� С;�4��Чjx��D��(8�GO��}[VJZ�(+�u�>�|�1 �{���,�nQk�Pz.˟�y�JVwMr48;o���5�_g���A�'�W�+���5�^3jz�M�ba��V�q�~d�+l�n��}WЯ�cSb���㪡73n�}}�)�~�����?�_6��m��y�����n"���b)�>��-5U<	��yd���Z��	��x+^���yб3rq��f�>�~�uD�軃�#�����PyFX�>m��|�@���5�E�IO5�%�v�]�.�F\C��j�u������fN�S̤e�Jp�f�Y}��zv��X�rӇ�����`F	a,i4vZ(Ui��G
:�yH��8�Թ��G�h5T�3�㴹����4��n����WWIK�+����>�sǣ��R�<r�FYeNBr��4Fd|��"�)���M�%�>���x.F��0��:BWXu����M��V�CE�>�_�����:1�g'�0]x��pa�N���R^�U<��'�6���{)%S�{�'�K`�V������|��aъUoWr����fO,�X��|aϼ �n021	ܾ�[�wBb����~z��J���"A� Z aR
k���JX���Q�s_^�}>�Dk�
�ݾb�\�`7[wj�%�4ݱ"��h�	MG���'�ݰ`�L[kD`C?�V��Z?�&�y3� {����\��?R=b�Q&�9��cB�Q�Q)#䷯�|1��ߦ��N[ LL�!WE`�"!�f@\8�|���S��;��+]&A�x��8�B;��`��y�|�<��<�&T�s�V���c����/P���| ��<�O�,��uw�#z���eM㫩5�hQ2�Y � ��w����l���sfR7���Zb��x�}�ԭ�_�9�������O���2�'	h4#�n�j�R��!y跜A�V��̸���p��0`C����]̝#Ӝ;V�*��k*љ;s�q�R0�FL�|m�=s�V[��;GK�H��8o�Vɯ� =p��K��*�M0wilm��Ї�^�,_֕�RI�o�Hzub�<΄�L3���6]ɼ7>���(�?X��Tu>_�Lc���n�$_��C����}�u��[�e ߒD��w��fX�Y�@3*'��b�c�ט{���0�Ye�X��*��I���ǊV�V�Fv���~��5ꛬ�y�����W�ZW��0�D�ksAq�!�s��#�VI��������iJ�J~Vyky�6Y� �M�V;l���I���H�}.�p 薠g�+���9��6�C^hO<WQ��y�e�6�}�E��濃�?g������k�a&�G�!�ᣛ��f	��}|�yn��G���л�q�'��*����~���yc�Hg[�(�P�5�
wV���{�ڦD@���W �a������/}���W�sx���h��U���)�����V���j�o��Y�%��{��1���Ί�FV>b�NWDk�˶䜍a�:*y����X��v6vԨN���P��L�ν��'�=�/���i����;b1�&�4U/9����D��_������)]|?��&�BO[7>����33��m$����=����f���-��m��.7 ��� ��Ӎ]`^�Ó��_I�z�&����2�����V�aa��.�K1@�|=�}"�~�k8��Q7U�></��Ī�p�{%G~x��c{��z=�3&�8(fq�:^~���a��ڮ�-i��T+0������M�[g���'�тe,��_������tS�QN��a�1���N�34?$���P~��)�X��K����+5�HK����2�>�_6��Nt�,D�z|�k|��h�
�{�+M)�K����:�.��G��S�?��(�hը��0U�<i�Î����Z	��w�	'(�˞68]o߫,K�$0 g�g��5g$�#�GwA� ��Wd�Ț| �\ϗ�t�ζ��]#W-�?��c���\�{��K~��?md�h��*������ᢠ�c߸8.������|t҅M����0"r�3�{9M���W	�������1�&v�pK�c�E�>1V�׹��>�z˚��t��%�âv���Բ�ğ1����׺��PT�|��!p�//�-v�U|����O2~��v�,n y�FUQ���q�I���%ݡ)@��m���?4���ޮ�V�����\v�*<�C߽x�j����z������V�<<��}F��ǽ��yz�O����4�⑅L4�MLڬ�[N�iG�:"��y[T;	���~�8��gmӼb/��)�;F�St�𔐍6�i�
_��qZ=�����:��'��a��J��*��q�qo���h�P�{T���:6/��~ś<��hX5^i�OԼ��+��.�',��mn� �0��^q)�M�p򇑊��*T�+2y�5 ju�v+پ��������޲�]����F,5�┴�C�}[M�H�-��Y�cV��(�r��\��bu$�C�6�p5`@�y�}G:_�!�x�G`	+�;���eho�d����W�I�i��*����zq��ݨ�֌�}H���=�) �����#�>� �݉^�Q�J��C��a�d(�:+3e8�d!X��o!�ŷ�#ˀ�I�a�ո̥�1�X�[��-;[Ml��hg�^<E�<[���s��r���:�R��C{^�b=8���:�V�˲D�6���S�w67���ܪ����ui�LG��'8����=1"�U$��I��@=��-��4��P9�_����Сa��LZL����o�nm)���z	#�����HXl�/�o}�P�{1E������vF��Y�'� �:��վ�qJ���������q�8O�k*�tx=�o/���~n�+���޿�H쓘B�Lu�nݤkb;$�*�� C�*d��.\i�}�±�[�<��"'{��;A{�'Ҵ���N�� ��kJ
������Yrp�]nٞ�>�DzH�����ć�£��F6ol�pt=�i��+g����Fdoh�j�.���{3`{��L���߲~��a��� m�i�+����Q�W܊C�f���}�����M�?n�я�,���|�1�#~SQ�p̻�����h3W�lN��_G"N���8:����\�6���iy(�.|0&�a�q�$`�{cA�I^��"��b�^�t#C)��(�E�vU��9�YZ����"a�-4���tW �X������)�BĒ	#Ґ A������SHR�Zc'��1�f��'A��n���7ݼ1b�6�v�#í��i��?�$khs�ιV�dg���hL�
`bn���V�-Y�3vN�jȣ�/{�P����c��x��-!R���a �@����ȭ."�� s��z��.��5O�7]+2�)g jRꛢ�۷Q<دt|����\=�������y���u��-:�p' �3�t�"�Ӥ��,���^�O(�I�
T��E��G�|����E��Y.X��c���p�SA]ݢ_�Fs�:y8�5~�*[u$������*9o���-��}��8X`��8:�<�c���M����8�}����M�;p�{���0�Yf�7Q�vc�;�R��>���g��N����OJ]��*���b�ɵLuW�{Ya�ىL�E�<�6e�66�	p���:|���"W��W�s �,������2�T�\�u�jI6��r� (^xt<�UFD��XkU�X��ό;�F�m���oǋ�����`;L�VCZ���Y��������j;���Iӧ�E�[&���0+*���G��u���V�fJ�#.�#�8��������k��'���b^Yq�@�Ԍ����|�G������S	6RYi!Cpu��w	��~�Vd)I��0#Ǌ�T�عz� 8���@T*������񄩎�Ǌo��eL�M�B���e����.�=3v7�aN",�!,`ڕr.���z�9���i�K �����1q�ނ�J��|ͮY������^N�)�9��Ocn[�}�ɤ�������z�=�w�Ί�_AV�K_D����P�U�|2���\~�\]��*�ӳ�I����~�"�'X���~����T�����>�I����Qw��,�v҅���*8�!.8V�P�<�����í�K�h�x&*SΔ~�{��H��9����[��v �t����Dc�������F9p����^zE�`��β���|�O�K��$��x����Kը���Sj��JDZU�>��{�2�	Y?-Tg
��`�W�0h�|v��$)�%12m�,�r%��&C+^/Ky�cJL�]0i�+�מ�O&r�+4�y	�R0���yT����9�?U>fS�i�MUU�����qt�������ONX�_R�N>
6Z� ߠ��)��S��m,���K�*�z�u�8A�-��;���N�sj�����%Q��"�b^p��o]�ԘB�o�� ���3B�]�����%������`�re�2�kG3�����|�D����7�����!u�WH�k�;{�p]���ӫ�~��de��v�s�EC�Q5ν�uC�e�?=~�?��4�V�l'�h�t:�pFA�fU����ܧ߷�6�F�w��À�l�Xk�Vw�lp3ɘ�V���n	����B������g�y�j���/�|�	��\�`�y�I�3��oV,<�I*����?v�t��Ol)��:�����,u�9y���]V� Jr�������7�U�)�����R��ؕg��ќK��Y�����2�[�������V�#��L��<0%'�,�
L�b�M��_�j�|^��X�ߩ%�/��d��yڱ�5q����4_��N&NЋh�1Kdu�.Zl��{t�1���9lL��a\gI��8"m"����qі2�0���u���4E���s�&�%�`#WJ�Vت
�^�{�x�0.��;���+�<$�UG1L��SK8��$S4"���-eD�اp��9��.̂<fAX�  �~����l��3������)D�ڦ��&���y�jsw[xM��9[�� ��"ކ��SG��6�NQ�'�Ң�f��3��w�	�Lz��2"��V��Ms�Z��~�S	K�A ��� ���7l�0#o֮#�����X/j+:�$�w��]�5䞢	��7c����6Z�lϏ?
~V�i�Q��[�0�ֹv����{$&1�⑲~ i��As�^�9zs����h�Y�#�o�{�������f6~6�s�aE��=;*���6�F����'b��I֬���.pD���b� �vOƷO���!�Z���	��=� E�f;�5���
�uȾ�!��R��<��0�w�[�;S�� �б<��w�e��x��K5�����y�S���N&��Ƞq�sG��$���_��5���k}�e���:�@s��ʝ����z��cDG����m �&�D ��L���I�_��^g��  �HA��~+▅����k�}�^ �z@5��u̍���<���{����)o7�:�9�@���?hZ5M����%%]��-Uƃ�7Z��;�g�=�3>x �j9�.���9&O�-��}���j˕3�g�4 ߈Dl�r���ʕ�ճK��6�T�e��R�D!���q��H\��w��J�<᳕�u4�~�o���f�BP�൪X�����)G�'���Ľă��K�.{�#m����,�P�B�X4�о'!��*H�R�j҆��u���o�|���W�7���So�C�~����T��7�E��iYE����__���Z'�l���=�DV��������uq�G��5R��'�sEqp��S����BO�D��o[���8!Y	"�}"�b_jp~SK~�]�EX@����K�m�_C\�6rx-f<�;j�
�'��I=jִk�23�|�OMv{9'��B�]�K)�+ÏQo�'O�e>��E=��ZxVqt���X������e�c��U��~h6j	�~"]��;��9#QML��)��<�*�z�O~�olSUNu��n�_�����i�n��/&}}��k��s���F�|,��\A+����p���{�y���j���h��f��Y�h�{�î�����7xK:�?"���q$_7����l)����]=����g��C�y��xr���Y�d҅�Q��F�ƾ�z�����o
yBkÝ�9ĉ̺���,
�"�-(|��W�����q�' ���+Q
�x	x��䃬�~h܎B}�`,YJR���g$g6Rʽ�
?�9��,x���]�c.���)3���ب2kS�!��4��B�,�2��9�p�{�уi9,�����4�1�12�� �v �@*ّ�Z(������=��a[��}����C눏I��}��T�&���![���4���{
���j�a~�IN���P$�����������͎����ӝUcJ{#C���8(3vY�I�n����Lu��ͯ�g�h��r_���Κ2���ڤ��a�!�([��fg���W`��G\��ٯ��N�jB��򣍟#�ke^u��	�!����i�BG�oe���_�$�1>�@�r��2�q� s����B���� �� �#�KY_;�;{��G�a���0/��lY��[�̸��}��ג|�+��9݊��GC��g[q�1�D�]���>�|=�9����p��.+���I�q(-0c%if��#}��蘾�@3�K�����!d'vu]	���[��(C>?�5GַȪ�9�\z6��
v=�	�?��˙;6Y$/(����U	�ց���G(�}� (�R�����RȤQ׺�Ab�����-�����u�Łq���0ʧ*gj#�'����7�`q�Cq����7H���s#M�� '�X�����}	�7־!��>��m1���8��A��r]��D�����}vù2�9]UU�RT!���/�pk5��:��w%�ʣ�>35 �yz��q����4�ܼ%T�>�qQ?02�5�y��������9K_��2�;�}���]V���<�A�}��~f�!�S��:���Sv�r�6��
�hahI�r�-p��a/?�<��vX�&K�:d��<+Ёx��Cv����f~�������lN@vҏ��<�m<�f���؁�х�������ͷ��DU��q�[T�R�V�S.A�q[��<�n.�s�N/[���,�܀�(�
x�ek���ٲ�+M�R`��v��5�F6ׇ�u��"���Ͱ����W��'���wL�F��Z�qpV��#1���˯��%zX�N��,lG=�㙋z��Մ=
*ψ�_����2N"�[�;�⮳?+����ç5h�@?�����M(!Q��e��XZl`�`�2	 ��|��zH���z!Fk9�'�:����kg�*��3�2���[�����p��^�Uy ��?����s�7��]X�� Yw�m��ſ�z�,��������֔�r��@}�s��@�|�����.T��z}�U{�s+f�a�𬴽�.J�֠ILV�WviR��)��C�Y���R��Fw.ۙE�>[�R����ɪ�_����xƑ����ekP�=ⳋ������rB`,�K�\Ru���'�Ń���ʕS&��8�
�Z���a%ʥT��ܶ�N�Wr�pszH˭����|(O�?	O��a2
�2�p �����˪�~�@D�η��App\��9�^8�FtìD���l����]h������
�WN����L��R��o��L}��|�to ��_�����r�=/�����d����y�
���w'
-؏8Wzf�Ǿ�踫������	�֣<͑X	��n=��Zaj�s�C�`ooF��>ד冼م����n��+�7aPB��aN"�7�!$�	n�b�Pd�T�#����ARI�o���$���8S2l����fM��;��UjG�hL��K8r�v��� swm���I����pZi�4B~p���4�A�/xf�������u����2�N>��j�e������Ԕ�o�M�u"�8Dh��2��XddS��UQ��5J��SӸS�9z�G2�y^�ih���bW�{pgK>���Z&��
Ж�lA��kn��k*��/Jdvrb�mdP|<o3�﯏��(Ѽ���/t��C�}y����W��l���[,��C�����G4��'I�����0	`ekSd�AԌ����	}+�)��ꡆ�r�Νr8O����[r�8�x�rUq��@�D����A���j�aU�̹�w:0��mf�Rh����̲m,�ذ���ܴk�I���!�L>�tL���щ�e\�8g���Vʂ~!L�A�ҹD�=s��%�Ef���(+~��E���~1�p�ݭ�<���b�||.L�'�:oN��A���u�����<��)��N�w���鞓��͒�����͵�d�ƈ8���D�.b��n-:�am'+qo����Vs%A>��ig 	h��)�2��'��F�J7E_ʓ$Ɇ���t��@���M�A�e�T�.����"��!K��$��qx�'d IXO�se�i�j�[0�o�����$���
�w�#f6M^n=�+��|[��b�ƥB�J�Gc��`���\6��O��W��) �E��h���L��J=�5�tǿ���z�&��AeC!D�@�����i��)��_в���ʊ�/�`$�:�5���� ���c���[�g��7^_pj���]���~�<���T�#����@ROq4�QWh�G��H�YF�xh����i�p�����O��*�I~/~�e�ctP��d�m�⦜�=���d�EZJTĨ�5Na�94A���S�����Ӂ~��
#�0���vD�V3hZ0���h���k7��Dz�4Kt&��`h��d�t��ʠIJ�@PY ���60p6���Σe1����'^�󎳿U �8͉S^�m<�gu���j�ɤ(5�������Y��
���%r4U�HԎT/o���(2�6�������A���j�����x�׿纶f�x�� ��\q��D�Jb�_�셭�k
{v�%��0���N�#�y�"�����Lq܍!�R��)>r"+C�S��Џ�j ��G�hͅ{Rx�����&1�ƾ9�
X�3�ޥ�m�URe�r�G#�$���v(�ZY�N�N��==/g��4uל����>t3�.��w=?h���e�p�Y<iZ�c8��,c�=	7�^.�@J������X6|iýDT�R�X���7/����������:.������,�eY]��;�2�ʷ��2.����I�9T�_O��n;{zmJ�����ZD�Y�b�A����G��o�������(54��q7c���Vt)�%m�����������E��V���V����_)m\u.#j{�`��=䴜�55�a�q����?K"_L״�8���ʂ�"@�^8�Iy��ΜpXn��*����L�����^^�{�c�y_:s_u�����Z��B��K�ӫ�Ym��!� �p�=o������^g`����"�Z�k��U�X:@���Red��#���J�aJ:�0n"]�Nbo��c~���-��a�XtC��@��[0�5�ʵ5
�;�$��Sv�C�Iu��R��#*(�A��/De�<\����jP����n��~����xGӢ����F���FF;����Px�=[8Ϣ�z�zHb�U�#·̕_S�X��fQ3o`-��ǁ�ͷґ����7&ݴ��D<d�++�ul�Y�͆-b�c�D�Y#_����\*�!�6�R5�?3J�e��ޘ�Z{s�еꫤi^�zs������ѵ��'�W��C��E"9����������������s�C����b�j\w�U�O��M����;��o)Z�-��{����	��{����%V��K�]��xPЩC�	I�ۜ��{bzv|v��v)G��KG�-^I�[��.������g�ݟ��SuJ���J�׬�.<�ֶ~��/������|=7����t�����,�u��8������`Q�.���d�z��x#����tQ��%}H�a7�fhл�~js E�6�@����⦒>���R���J�7�vT����]xIf�UX�Z�s���B����:�����õ�=�HjN�P�Ú�a�����#�9�{�/A���̙;���9&���ڋΘb��L���1<]�)��W��J�c"�:�+8Ď��{4�#�]��umo�W���V)N}^
t������<Ty��N�8P9H�e�7�)�����hhLu��*Llz����F��ҧ�uVo��uS��Yڪ�嗿W�I��b�w+'����8�U�Un'��#�đ������vHhT
�5
l�Ζ���}T�z��(���t�A�0��:��ϋ/����vJ�6^�m�y� ��ޝ�6z*{2?h�HQ���E���&�������a>GǇ�8Zu�J�%Xu��\ԣ��x��˘u�@|���x4�}�>��qkā!�7h+l��BT��#���`@-�ga�����U_{����3��vw[74a�ӿB�XY��ёK�˱��G���<���=�k���.wWذw�O��wno�Dq�[}�lr~���e�>�/��>5�.}jܿN[.�� >��c�}V��Ìᮯ�eps^�k[ȠT�d���4ml�O����m�-�vL������*���������N�n)�G�j�O��J�+�d���B&�^�.��loy�9=ƇI��i��f���W�"
����#Ńȸ�'��c0_��00��qNsb�L�cW#|�����ʢX2�ޣD�"ާ�qA�$�3,zj���[�n�E,
��Y�>ͭ��|�;����[u�2i���$�֙f���R�R��П]�w�kd�.��ղF�Y=�g����4��-1�'#�D�=sc��'?O!>�$fV=�I8*B9��<��w|���t#oܦ�s�T92�}�/t,��ˇ��;�}O`�F���|~u�[`���]_�ZB-iiބ�����?�L��<B�Cl��e9"V�2�U�\F;�bz�	(?
�e�Q�+Q�=M#�Z�'������O��9�*}�h�ӄ�������F�Π˱�vԚp�s��UŐ�2S�����t�J�]��J��0ťv�c�rM��a�.��uWsb�5���y�؂� ��xt�h��P����x͵Rڠ�oeї46�M�J�_AI�a�̠����R�uFVyP��S��DZ���şhV��}_��l�1`qZ�F��O��".�_&��0����9.3���а�[X��1���a��o���x�<`w�r��z�DC�]���vp���YB����x�����g�m�ȪXm�6B���a|��a��&�Q�8�G2Q�r��L�(- _D���净�ʂ�&<S�l���*4d[�[����fW��:��l��o惊Qa��Sˎ����������J��A�4S�O�G]O+#���� f�ǃDѨw^��D��/)Q��GM�����̗ mD�͟ǆ?�H�d����\Y�+֒2���nB�M��o+��۵������3n������K�S*�t�4�q8�r�g	��迫�_���pM)IRE̪��';e��/Zb~���_���?c�LOM�ㆉqN7cb:�M7��4ӛ:����Sӱ�s�4�tǏ}����_x����~�wRT����9�dl߹�E-$��J�`��P3\6M���
��<HrQV�������!�oݣcϋh
UT�!S�N�7���]&������VpAYB�K���nU����XM3vц����b�_e�35��|4�*���O�V���+y%{�A���UHYv'�Rj��������%����ؖ�����Lx|y1p��0m�25�>ލ�%�����\ �[�+H"y��C��l$�?�p��<��@��sx��"��x1�Z�r����De�b�r�.�.�W��"��t�z첡+��Y7��T�ћ�E f�)6���ėH<_P�W����gI���80�i���0�Yq�!)z�,R�]g�řc9�z���K��~>`��VP�>]#)
9hM^W;�<�i[�I��Y���]u\�z��$�c��i�7]��h��K�7��Z�t�Ji�|��#��y��sN��YJ�Y���$B�S�����}P��Vғ�;�'����ir]���Ga- ��0�}'���H�\t���Ɓ�.��l��O�Tu��".���sL��?�}~�$�$!د$z.p�
��챍_���2K{r�R��&�Z�a��J(WW��>OYQ��5z��|^�6p���Jq��!�R�$����a$R{�W�(/P}:��wv���J���CYx�X��םcIxdf/p��]A�'�6�h���&��b����(�ln^7�*�-��xþl�n �"@�/
��>@�o��=�K�X`��� ~�km�8�JLu�wbT��Cȣ0��fY?�����Qw��?��Dx.�u/�nwj�ҫZ�I҉�!��g��QN�'����}q����׸O���S��J�˹{��K�Ī(�M���zn\��y��y�.����l,�0���%f����vM�t��z�����b��T���r7�ڛe~�*he�{��)=����,vU�4�����OO�Tl�je\�gk(̥@O�Bov��xCOV�o�Ӯ�]qx���<�3��0���i��������
r�t�xM�kc�kᤜ�g�ޛM2����"w�Kb�t+�4U���q���K�Ø���Ģ������&hةC����_��F�°�N��Ӊ�+78����V���O���Hu�(�6���%p:7s&%�z���Ǫ4^��ˣ�6��mk�$.ƃ3���L� q��3��D6L\r
{f������>��
Z��h�|׊�E˱��5k�A���	�<BZ��h�L��;�]��K_y�*.��|Q�I)�p�MVA]���>m�V!��\�'_��>eܟт�I�F��Y}�[Nع�aDFf�^�>�"�dG-����Μ_Ћ���k o��GyY?F:����͓x@���8\�RZ��W&�^��.:��M$��;z�G��;}!��9��`x��V݁� h���#�?�3��~I�h�-��!9~�h� �G��фFy$��,2�V	�>��$dI�!��]�$b�/ ���G��� c7�z���%I�77Pt%m� �=O:.�.S��f)��̒%�5_v;'b���W�)�l�K��髲�I�MK5+6��m�ف��'�I���\�C�b2�A���������>���j&a��s<�3x�֦��Nk옻��je4��i����� �m�w¥uQm����3��êJ}54��L���X�Xy�(`�s���MFNÂw�-�Ol�F�M��[�C��ϛ��͎�ˣ���`����ѐ�GnFj4˛XN?��e�y@��Y8�|���p�O�?I�y�tӄ\�Qb�s<�p���؍�,ި���9�7v�n�P�5u�m%���� (>ܘ�'����S2�&$~_~DAUiA����`�w-Ó(E�y�m�ؖ��4�:純��>iw�;��g��g�Sw�j��fG�Hz��+�ʮ�~ip`�%�U"n3x�]H˷b��k����f���>��6�Wa�_СW�C;��r	P`Т5`X��>���on�&��c���c�ĭ�'�^���0�o�����N�`�\�:�?��:x���7�����o�����[We�������:G��pЯj_�J� �!]oӋ�~d��+�b`����5�K� vV�1�.�G��J鿇()9�~��	�<��	��9�x��~�>ۍ�gS�/@���5��*hҪ��@.*��1E4M���Y��G���m';��Y�\����o�Qr'�"��u���att�O�ë~ۼ{�w�W#����D�-��s�H�)Lx��k^������mc���{gG������Q�Vb�����/�a�e8��u���(��̄�_w�7cyc��e�vL�֥�9���}���tN"�_�pJ��|.ӫ*�/i�Q��H:Q�9	���8�$و����F�L�xFhKS�6t6uN:ł�t�,"{Ya�B$o�ӹ��P6��ܟz�m����B�w���Q��K� �+�Zx�4��jQʤ
.�?�I���t�s�m]Ap\ W9�����j�Mdpy�m�����S/�<�\Xw�ﰷ�͚nl�����sjd	N���_��WV��*��ʩ�@��%���?������G;�|�Q#6�:���Z���Τ�����(�h�؍t�����δ�DA�]��Fw�oğN�+��b�CX� �ڛ��^�N�E��ZB���3~f�r��
G
�/w��5�&�r�*9Sh�>8�J*�glTD��#tE�1I����/�xF����~r��ݒnT�y"�>���}y���$��d�v�M7�_���� 	]�M7��7k=�ZD����� �|����]!t�����m̚�d���ِ;�E�Bұ�eK�B�1G�$�w��6�������mL2�2D��ra->D�cߖ��;�7 �T7B)���+�ޏ�v���!�*�3�{����&�!��*��ܬ?N�Ĳ�pyx+C2�������%1w�^��Q��6H�������2�=&��2��:l A4�u����W���C�#>n�Y�|��9o���l�Y��yi�������
	WV]�r����5$��r�w9�+���|<Z�����N1��my`���i�٩� !�27̤�7l�-�N�����}N=ï�g6�vI�&�_4e�������N.�U��]��=���͂}(|l7h��L�+��T����O��f���0�(�~��ON���h����F�b��ژ,U
��@G`Y�� 8)� ����<��A2j��C:7a��|D�+��Væ����̏\	�R���(R�q��\�q���]��
�Go��#��L����57��OOǣ��d(�Vק��/�[.��9W��.�W�&��)j�<�r�"w~X��M���A��
��x�4[�s>dj�3��Ƽ���׽҅ؼ������n̺<J�
n?���U��S'�����Vn����w/5�Lӈf2*�Ǉɰ�,�`:t����i�0o���^.
 캢Bq��ďn��..����;(��������wh|��H���~wd�f$��7���O�Kk�QB�[<�\|���.g�ꃟM���R�g,� �I��?��M��1�O0V5�>�dof���Z��v]��9���gl���tE[HNn�I��(�כ)�~ۡQ@ϫ��#	�>p�O��5�؃�����淯}��d.��j�V���� �09B�V0;���(_�L��5D=l�����N~9��Df��|�� ��t�9�6,A�N�D'r��.�����o7�S�H�x�G"���=������~\~sԣ���U>��2l����sB�π[x���ZC��GĮ�~ӫ�%zҘ��H4L��i�����X	vgN�y���	0��~Gw��^3v(Ѵ�K$�~2ewJbB��=A����|u�w[wl|	6��~�f�7% �KC>M��x�"de<˭���D�@G7*,&�3��9Kj�!](��ܞ*��_�K��}0�\���⦟	�����r� �E���m��_V۳({+�� 14��>�^N��d���S;��\�v�I����������o�<�u�r��Y��i��Tn�LمsW�CD�eS�R�e����O��*xL��W�jq:|���A�_9X��+W�#�W��bY[(��M��Lb��ܮs�(C��?�֞�JS��/Xz�)�g�����s�U{�%�͜w\��i̐$�� G��r?wԮ���~ʆ��m����8���|{ϣ���+�`�[�=,���M�]i8[�,7�)��BР�|5�Ju :�#������JS�N;~E�|b�wz�K�B���׹��������T[GI/�6�Dv��%fB$5�NJ��!�,2�ğ� 'ZV�Hd�қ�ĩ�S�A��2�eH���ro-��L�_3.(�ߊ ����UBBw��?���`�W�Y�գ!k��G�����F�v��MS�|��8䘾���o�`u����ˮXI�8�ޕ5an��E����E�'l�$�7��Z�3�'�����b���HO'��~R�����I�ք�H���Q5e���a��]�HV�O=\_߿�I~A8;�g�W��A2'�'3�L?�-�[�J��W�"��&���-�l��xث��IA�IL}��c��R�E|̟.=��H�J�CH�����Bw����Β�c�"�Ѱ�޴D��1�ݕ�K����;뱇^���Eu�UW�/6�⬝��.�J���Zbcc��/�2$a��b�+'�ώ���S5�L�6�z�tAk��v1�O"��g�f�}����v��bF�]ͷ��8^��@K�^�~�����#k=MfD�wY�	�au��8�z	~���yY��z,.�?��۔�l�ܕ��8~_w�ȉ!,�ig�z���1�JCJv,��v1���E�}SO�_�*�
�lV�L�x��4wq��&�JZ	�I]���q/�*<lTB����M�m�q �H��I��/se�|�>�����Ӑl��A�Ⱦ���s�x��:���+�mpE�����2U� \���h���p�_���F�ϔ��3��]�=��d�Z��0�
��8��ڧf��6��x$A"vk_ۿ1g�/��^6耀�󏹒�p�p��̫���lq���V-ffW�d���y���O�%���D�>_O  �9s���졞
gȹIෑ����N�x`O�K���C�;��� -�tt�Ӧ�'J����U�t�6� |t ���&_�T���R}���}%{B��&N�dWR�<���{'zi���T�F?n�St!li��@7�+W��=�La!��H�q�~r�&�tve���F����^e@A�r`�Tv}8ofccC��hu_�arӌ�T:��]���<����F�j��7�^vb��>0򫺤��u����[Uӧ��?<�8�5�(���e�aȲV(O�eD�$��l��pH��Ȍ� �ݦf)����]��ͳ�Y׍	W�4r��������-�38������֮�[G\�8�Q��ܜU�s��)J��"ck^��7-�Y�����Q\��v]zvr~�����J��]����������)��.+�v��BZ�?J����e)(�켠ϲE�f�[�A��o
�	Њ���v�/s_5�������j�w�s`ƞz�F����FLg�.tR������s���0���cGkx��>@Y�IH�MO��j�O1txg�y.H�
^ ��%��D�v�;<�_��f�E�9�7�����;b�9i��,���#vӁϣv�=r����
�H޼�%���n0�3U�&����_R���&My�C<[���"�>�^9/	2u�ۛd�.hZ�f��P����:B0+��O~!�P����[q0�N���Ϝ�+/3:�4�f�)�=��5{��S�w�^��q����_s�Y��H��hl��~��^H�ea3�&|��_58-<n� 6�b�>��j[z�v -G�/؝������p��Ty��?i�?�Vt~�#�pE}.ʚw#���׿��ͷ2��]X���c�_�!��ݝ�e�ؓ��-&Qe{%I	��}H��&ׅ��������جDc��?@�?C����f�KB��������zj�&������Y�������՜TF�,�7R߻� �8�D�H�#G�Tr>�M-yQ��p�۫��'��,��}����d�����T���t�|��*�4�1�h��s��m�/�Ea�!L�&���)b̜ eٓk%�".=��]'�>j��m���7��	Q:�����G!U�Ƶ���_8�=H���l��m5�#1����2��\������G#�{M��i��O-`��A,��M}𒼽��]9�����5#�Z겳
�������[@"�Wc��+/fP �a>���'���KY��A�}��T�EA8�h�d%Y�-�$q:U��a�]|&<j�R� '���LR���:��L�J7��b�Z����5V�V�����P���y���n���o�VN(YV�$
`nz��}j���ף�F����1����V6�,o6�媋guK��~7�VG�bc�Or�*�=Q������{v�+Oݪt؍�w6��y��Z/74��h��B���:�/m�d@��e� �C/Y��.���bS�]S~��?ܻ�$Fh�H*��F��`�SX�F�	��N���
��,{�`5/_$1�v�,7�P����}=�}ѕ�-br�M�c�9d|��1��s#��3�4�o�Q�z�5��SRd�}�&�Ë���J���OW$'����h�5�]'�ך6�Ol��L*�/ة�Ȉ\'3� i! ���ú�5o�3��h���r�Tm�}xx�`�+��5���S���⃊�{׃ۿ����>sT�7��D��$^��CO���?eY�x�e�����+�^�viO%�Q�J�1���-a�\�2�H���k@iPCq-�mt��K?�'��;������ r���_SY$�Y'5sl�R��2�-����TU-�*�Xp<`Z��oHI��u5w'F�h\��;P��һ3��f0�-��=R޵C�A��XR>	�gʖ�L�Q�����w\�W�U�L�C��dL_K��]�C���oDQ2��
�`]o?��o%Q*Q�7$j����[T����07{�r_��mc�V#�Pt���p�������+��j�3@�L�����1;t��!�j�wK���h������
f�{�g�\b�;=��VZ0�'��x��J8[�����+ˡlN:�q�n�Σ�J4]ι��)U�w�3�q������� jP���(}�~3�V;����Aـ2v�16������Oؓ�_z��;�V��j�J�9~��6��P~6��2��c6������.p���A+İ�ʭ�Ū�W�L��z6�O+x_T��bE|��2�X�#�0|� P�����)�CrKv����0*�~߫���B��� �ΘV�yyȕ�ƴG7���nD�w���H���iZำl�I6��3���@]��v�5���,�^�<���v�h�������hZ����n馊�=�݈?��"����2�~���aCfP7�O�9S(~�g[��_N�a��ݏ�������Z�]��0���GphK-�]��P1�O-O�����L��N������i8�cx��V���zAg�ϝ�s�=��f=o���Գ�خ�A��꦳"V?K���ߦ��s���g�շ�w٨�*ַ�;��a�M4a��cT*\���2�$�&��z�\& 7�f�v,S����ܟ���5�0� �sV����i�� �����n�f��i��d�4�V�V�ܞ"
�F���� �)�Dfݨ��A,�5����E�;
%I��Ш���I�~��N�"-����t�aF�f�$��P?�I���3��~��Aq�IW�m0Y_B���[R�3;�1��z[��=Z�΢U��n��>��\���m���f���^�_�z��5,W;�C&1�dΡh#��uJ�z�둥na������m2M�̭Ϟ6�z��tRIE5����D9Z�u�(NU�6
��%��|������@E����0��;�����!`b�|K��y�3���ɦ����m�Q��鯇_Ed;jS1h�oFqSHX. ����l��p��"�zu*�)Fmh�V�7��w��;Py�I~���c���z:�p<��_X����W�B<oYd���Ȁ�Y$�˩�Gͨ�r�}~Q�G�-͛��T 1�L؁���Ζ��w��;�cYu�]'Kz��!��xu���!�Qb'*vrgN^۵�Ñ��~O
,C�(�֗�S�Θ����f�Fɍ
z�8f�/Y�(V��(����md�V�I�㛋����ab�"w��^��IHKkW���T�wE�6:��_��Z��$˃�T����3���1/�3/�5Z|Q�=�߃�����,>RV9�6�� $.VA)o�F,ˮ|n�+<`�V������WSB��Qng,S=��+1~^m�2c�I؋e靤�v�O93�'��_բ!ȟ��=���^����,��Fx��t�6,h���[7�#��e��%_)3����+o*�8�2� ;1\�����U�D�*��QD)N�c�t�rx���8^�.�>�`���a�@o#�x�\]��Y��p�Yt��[C�s��~M�[̽����ƍ���>�t�Vt���b��^1����%�O:��a��r�#���	+�uv�{��! R�c75�o�,?st��a)�N~��B2-�r��Ȱ�l��w���-�ȗsY��PD
}�mp���ل[KܯD���a���w�������e�H��
	�[l�>��ڹ����g��������UCL�W�pv�)���2�Te6��)�N[���4
���vԆ
�u׵�L��7%$~��Y!-e����4�f�4�UuLEJ���?�ʟu�qZ�Տa�iA�����;H�o~5���c�Ы,ce?���d������]�y����]����aR#��J�W�b�'(��tI���2���g�@Xk��a<?N�Ea��Z��{D)m����Ga�5/]�T��Q�����ۦ��w�{�vի��pE��5�dPY��s�r���/a
� 1�3뗰R�˧t����Ժ�w��Ux�c R�t%��XB�k��wƔp�(՗lFﶜt9�vQ�T9�Y����IXO���N|nbˢ��I+U��3��ڎ;H���	]�r=�:!ߏ�zc�ܶ�&YJ��Ʌ�/��|/\t�z�ͥ+���?���1./O	/��߫�7�[ޏ�r����Nv�w���<�?bCz� 0�{oAKC3�p��3���0���G�t������5C�- �����q�yv@u�������e�[j�)�Z,�#jJ�����46	V�wGྸ�';ϫk%��1��pb�}���mji�}��TY�����#��S���M`(N�8�'Z�"�5	���<۠�b�}<&��1��̨Է;�����t����j�#��ËY��H��k|���;�~Z��z�����c~-|������/�4����Q,%����G
J��!>=[EݞDv�D�DKF/2�٧��"�CQ�������~��wo���"�V��F��|N�Ոd����HH���i��������Š��������w��mߊ��HR?Xs�l����}\*m8TƜ��,��fݝ1|=�(�TO��P�j��&3���wR��~���)	2��z��I��b㫫o�h*y����3�ΗL!_�xn?�ay%����4�������`�Nq/�H>V�-�hĎr�#׹:~�8�@�!R?��8Q�]'����O[\Ij�z�\ϛػ=J2�򬝐�M��IW��j��㸲��"�|�ȉ�r�W���z>y'�HU ��,</s��+f�ˡ7����3� ����ޑ�a�g�mW�ID�au�rbەrgp��5t�& �n���ҿ��	J!a���O%���W��པ#���slKig�eP�ү�����i,}�Q�3'�x���@h�}9�^1*B�(GC<�A�^2����ue�t���� �$L�]u7؍-�����yZY\�p�d�Z�zLĀ���H���E�q�V�X�z\k%0�����wt*���$l�Hǎm����j��#�t�E
m�5t*�rm�i�4���ʃԬ	�&���v���Y
^ЧW7N�[�	+{p{���/�^�\�[^��w���~��Q��p� ��}PO�hÂ/���x響�y5�S�hh���)�02+���c���s�\���ơWx�}��Z*�.�*��\��M
ߝ��MS�4��r���.U2kE�-0�a̪ZB�o�ܮA���:�$�vP���O��=u�|��r��4�dM�I��zN�hO�g����Gǩ�S��m�j��b=�����c�[��º=bS�{�(�����4��uW����'�G_��g��÷�ZY$�'�*W��U����·������6:�/￟�lA�w���?��u�ϕ�}Wyii2rA:~�ϝ��Lc�#��%2uh����έ�?b�c�R�g/u(�����I��¡�xF��������G��#�wi�H��7�iU���`,9j���V��r@�_�$�{�{���2o�tVDJ��Ͽ�SJJ�� �`h$T��g%WMl3��湦�(,/n������V5'�;�9���WJO`k+,� �Nx3_��6VvG�9���N�n*�B��ׅ+���5E	�]"{��k_���"�>;U���;�ܪr�����tDMM�{r�z�L得G?P�>긽
%��vCo_?9�{'���yZ���u�	_H�������ɩb����X������-�dˆSB|Y_Ԓ<����g��S�,!�x�M	�*��+�>��K�3V���c�f|���gy ��2B�m*���U\I�L��(��o��#��Z�a�6�3���>b��g�|�+�J{�*t�S�֨�.���S��Ԟ��@(E mMs��hnϿ�>U:þ��K����wUp��:ɭbG1U���Ak�D��ۣ`���:6Z����K�^���䒹7���0nkѠ����\�׈����?��������w[��#U��z�1����h�p{?�=<�rs|�0��.�ŀ=3���a����1f`���o\v6��O8h�R����E� �G|8x�}�ΗYHJv��~�.9��w!�;���?Ҟ6v�f�d�����L3�o�����#���0��B�{�w�ʲ3�U����؜��/Ͽ�"G�zLJ�΅�ʶ}�e&cg�ָa��'�l����E�>����9���Ս����B��!u�?]�|��P$����U��b�Nm�+_۵,�n=���<c�B��<RW4�k�
�v�Dsy4H��g_���ߞ�ڀ�G���򴍼���{Q���3���;�-�H������KWYi��?��h����|��Q�^J�&�em���,���^v�r)���:��:C�b
�3��,p�nJ����/r�n�gO�zqɐ2�Z��S�)�Bcv���J�J����!��t��K����昖�+�\E��2�_�wr�J^ś5��fN!�LIb�fF�;�ٲ��M~nX�>�Gr:��K�B���Kg&'��#F�;���2�7�=D*�&?G��2�מ�x���$��).��WlyZ���p�N5��M�7ay�����Z������^��kr�|LD�������J�q�����/�Iu����H�L��E�-����{��X��(Rq�Y�şM�L�w�8�n�ܨqU�R*1�.M��ȩ6%��X�s�Ѣ9��O�����8�I[�3>5ᬎQwh`\ݟ��)1�$�g
�.�S��X�T*ޟ��C��:���3���w/%1����Cy�vhB�ٯ���j����N�ke�k��˺������̹�?Ƴ�뱶7���r��m����W��Qzm;?��;H+\>�t�[��α���CZ9Ky�F����
��<�}:�f"#���?��K����b�{�ҿ���R�U]ޫ������k.�F��P��I.*��::0�Nf�����2����d��b�f���F���	˖9�{����R���?cDhR١���,�Q�w�߯x-����2=�.�P�}�/��<�'E��� {1~`�R��ei'�fq�M�k�k�#+�� {�o��e���I$$�lw�7�`�<��]&t�i㩺�) ă��ɜT�|�>��,q��v����껿�ک�V�fx��[��:bb�!~�N���I���H� �����N�����=/�Vl���*|j���YK�S��~����`R��'ȹJ���K�sC�n�mos�;���������������{�g���m���_�/��_���[ٲK������!����?җM��ʓg�S�ZVx�Z��Zls�t����	��[�Q�P�
�%Q�D�9���<��I��9�v�Ms^���P�9j��~�ߺ����k̅�+�R�g����&�5�9G>\I�n�ZuS7���-|w8���js�I޹ۯM�>3#���{���2��*������KУ�ck���[/Y����Oٝ��ҽ5_�ܷ�*�y���H<ho�a�$�b�̿֠g�����ۚ_`z���r�G�wn����vy���n��dFrr�����Ea�AK��_�������	����� 7�s:Lٝ��_�K�!3���e�i/��d���7i\�o,R�	�~R�1�Fr"�=��͠�_�Дz���:"���sI �&�*ek^�b�Kn\�$M]=�:��4��M��Z�0��o�,l "!�c�}8�HRs��[�Ȟ�+����З��B��
ڈ��ō+O��۫s�m!�~/�7��P?�j��5��[�����������E����o`�6Qyzq��B��g*�ܖ���-l	-����1���F�·���2��d˅E�o���Ԁ��T7'TA���r��d�WI�i	�--���q{
A�ܳM�)>��8�I�.�����=�x��ӝ�h@$o.�|=\��O[ړ��ߛ^ܔ_sE8���'C�K�ll7�~�$�^ר,�E[ד�*)?s@����ZX��t���9�+��[i^�J{t^�|(s�����#
�W8˘�׆b��)�Q4��z8z�؉����`�������'i�Ϫ�_n����u��:�=+� ������5q�lYx$&[��ĉ��[7;�w�6�����E����������2��'L�x�#��b��kQ���nS���N��cs/N��~��2�Vsp��=
�BC]з��O>�gx$��Y}F�G��K\}r�1+�t�VI�t�/1#�һE��D��gi�6��~�4�� U������w/+g��O��ދc�'>�b��jX�9���v��D|������D�+�^~���)[$�V#��*���p��ŦI����� �Ԟ���&;.��@��ߋ�_x�Q��[V���W���z����x3�����R�W�;�u�q�7�f��[MEs����@#o��n���0~ �e�V��f��DGm�^©�Va,s{c�-{�x7�Ӆ������6��W݅�%`�Y�9?*\���7Y}��\��;�9���S[`!�V_�0/T�Q�"ɘ�p;3b��z�q�c�H�Z��p2����ˠ<�Z�Q�D�^D`J�4��ąL�~4J۝{��g��Ň�?��[x ?�
�f�L썍$6��߱`�!�/VD��	���Ь��b�1y�*�d�D�x��w3�Ϙx��X�����G�3�N�G8��Y����� ��,:��d�8R}n�c;�6E�>��.Y�$a�r���y�I¹5�f}Mm7{r�+rN���I/D�g*��3=K��>�Zu.-��h�q�Aη����S�.����� �STܡm���I��4ƜT�7���!��n�=���~��m��� QT���IɈ����}��zX�[��~0��GN64mBb��%]���˼�������Fa�0#���A�P�VW͊���{�-繦��Ƨ�y��$B���"�ɇ�ؓ(�?���=���TϤ��,���utH-�y/���Wa�h��-����Y7w\��Yozض��am��:d�]7��iP�=n}*"Qm�s�ǳ)���Gi��U"���E��b�S[+�%����;�d�`�]+bǔ�3gz�����s<����Q���w~���g�nd�Ϟ4���H�Z��.N෣��B�s-����^zD=.;
�^�}���SS/��x����n��kie�gCvDe�Дƺc��-�LτG��H���BI�ߛo�-����y�A=�|�����fC�?,���O����hʼ;�n@T�4a�Qd��_938v;�yx�.���,�<��2 �*��g���(Fxj60[�*��9�[��ilʓ�*�p�ͼ�RMo�=�Պg����N ��(�Q��)V�R�!��c���Dm޹��a����?UW�x2�S/Wwu1��2Յ���-*$ �G�n�-܄����Ġ��j�^>{R�d��I�\ڻ��K$n�瑡p���c�OA³B��Z,E�D���.�Ԭ^@F~�R-�ǵ���.]�v��&c��(����D`��d��z�9L	O�6��s1ҵ�s*)Au�)�F�f0�$߅�Y"Xf� ����t���R�N��Rh��T�8�]>)6D��p��p5�<X��\q�L���o�5�a�0e9�5�-���V�oV��
����[�qG��[�)S]V��QD5������i7��Z-��z�	������v#�S��b����MH�G)��u�U݄����4G;Ԋ���{C���u������⎦9�y��t?1j��9D5�]�93q�(����o�1T&^&oY�����>%�067�������� �e/k�F*�jT�&�q�{ϰ>E�AGTf� Vr��N�A����Y���JG��z(B�	�IX\F����20ũFw��wz:���w�*�yҿn�7V�I�!��=����d��Ī��"��k�ݯ�N����>�ʖ̨�_l�y�,Dy-�a���%#�^�*?�i�c���-
��^]�kMF��
1P�����������?��9�TM�ňp�׭����S���'������������`֞j�����p�jV[ĝ��.��y�5`�������'�i� �H &r>���R��K��S�-�(,������ ��-��uGȆ޽g�Lu�Ͳ�Q��WP�[?�s*/��R�}������3׉�y��-3c�e۩n������z��7L�)�O�Z��6��/.����_��&w;&����E��?�{N���Հsr��_�Q���}v!��[@>L��🈩�����y�c���&�0���3_��O)}��I�_kͥ��+uX�ۢ�O���Q'�V#c3��o�
~��:Q{�Y�`7G�X�s��й���b����4���� 6VY��S���W6�,�/��.�^�~.,>8�>$��*K{��+
��1m�M�?2��=�-�B�Eq�z�pY��6�W���wBƓG=��n�����5 tq
[��Lh1����	6��L��?�"����Y/��0�q�C'�R�|2��#^d1x"qu�-�S[5�ݱ����k�,e`uq����"��7>.*X��n��zD�~�	�ъ����狱�(F�]�*9�{/-^��c���"m6�m��6]��R��z���
�����<H�W�Z9���ǵ��e���V4.?i���8��Q��y��c���t�\�rʝ)�*L3"��9�:Ed�e˝�7�B6��%��iH��bGO�UA�7^cuƶs��py�z=֥M浵T�����'���(�(|�u
k�'�Ҹw�Щ]-��UX.Dt�.�7�Y��/l�$j���j7��6�fx'>1�����������{ӓo��.���-hƺ��g�EvP-~Y���|��(<�e݉��n�?��u��?�M�Ŝ8����ܘ=����t����'8?��QXC�z���HF�邘�>�q�~��.N�8G�e׿r��y"�/{IH�}��C&�X.z�kK�֣�`��Ja�"�|'�/�H5����+g�Ώ✆9��ȭ��ޤ�#io�n�%h�����6��)ZS�-��)�ђ�O{���wIF��]�C\�G[��wӎ�sD����bh�G*����y�d�������Z�Q���U"l7����]Ե�gag�a��փh���3_��]���-Z�d�(�G:{̚o{
��и�M%�@m�v�ӟ�=�63R>D�98�[�\
of٣�F�5�+���8@��*@'D�v���G�����zEZ�-�N_f���T�ZP��*�#����5;;�&��޼6�݀�[&��`��;�bD{؞:\F����X�~;,�*���~�����q'J�$ҳ�f����F�>` ޗ�[����?��ß����$n!d�"��.)3#�쬬�M��VC*#3deӵ��h�{��{��{�܋k��}����y��:���}>¯�7�Q[�3����j���f�U��.�i��p�����5.@y�S�݅f��V6n��c.���qd�h2X/&�hZ�\�lu\��W���?���y0u��_���ͻ�^�x]�~}�J�Z�7�g!�s�ܵ)fJ��R���uP��\vI����L>Y��|��B�ι�:���	��p�K���T�;��R��\1&��O�U)c&�/�o#�#[ �l��>�����F<�ؒ�P�/7o㶎��*�O����C~\��o�a��
�|ٙYFܫ�9����Ceբ��8�1ԯ�����[�ܬ��-^�2|�1#��'!�ۅyQ���J�Y_�����{ێ�%wb;��)~%uF$�����,� O<��H?�N��v?NP���>�~([�����2��?��S��:����+}-ÑZ�����\�ˁ��c�1k��:��\��3���<v���HDa1�d�%j��b��JED �{��,P?��!%(#���qN�ؐ~�?�2zov����Nˈ�t�9�C.H�M
H4j���0Ж��7"�f��*>p�IQ�ش�rgR��y������jO�4*t��G��	*g<ا��,��)�M�#�+���m���U�r�ն^A�V�Q���-x�}~�]������j�4J��K3rrìF.��Q�rNC�&tu��E6��$mI�ξ5Ŕ�tf�$z��K��%�8-�t��uvH;�ؘ��j������˂r��ޓ���*)�K%W���:���ztH��r��K ��ߵ���h������ٖ�K��F,�d��7�Z�?u,|t/=[2a���Q�GD˃�=O.��?#�3U�E,7W;�����{ľ5Z�AI3�h]��<�$����T����rG{Ky���,�&aB]zy�U(�子�JA5����Rs�1�9�@U��:��ވ�6��x�N�X֩6^$�bXi�|!�%�=�i�����Wy܂b-�%�3��g+WT��!��z��oU�(�>�Y�\�����;�T�����\1���4n	9y��(��l�����js�CH~R	���/6���Ӳ���\[��Mi��ZW����C�~y|z��|�m�y1�z�w�\�&6b�1�&y`d^���%���/����5��6�~�W�3��@��`����h�%VY᣾d��=?�YI.:�wl{> W3�D�y�rN$eD���~��M�
�޾���z�p����f��`��� ����&�xk�kD@�_A8[�b����"J�����͹��>���*:��ʓ'jd�������$���ݕ ��;fS��y|K\���s�)y�6h/1�� ��Ï��*�N�5fd�g`�h�>I�x�[e�K]�S(*c�)���w��:Z����[�h,�o����=����׮d���p��8�Vj h4|��L�� =ZXL_Is/r��~.	�^�b�-J���B���^�b(��.j^�FC7���������@������)#r�w)oM�5*l~���ʍo2�FTw�
�f�iv�TS�J��	1��T^��
2'3M몀�o��+��h�(�l��Ƴ��j�ڷ$L�r��__�]k�n�K<0)�n|�Y~�	к�a��Rz�[&�$吒�V��2G�{�w3;�7�����3a��a�1���;z
�'�C^UH�^���EAQ-G��r�X{�}����MZ繄ɾG����[N�N�'Z���/z��?H�5��}��\��
�K�t�������ޠ��?5�T�=�q��fQT�����x��6����a�Y�Z�cǸ��a��B�TLL��n8-#��=	�N�����)���K���2�ۗ��f��)��+�=��'����h�'.dPo|��)��-�׀ �x��$�D�$��Aޅ�G3��ǿԺ!4�c��I=��d� �8�H���<;�?�"Ec�&3*�ձ�^Lf�1f�k�-�<͸�=��x�:�W/T>�_��X-}�|z�-t�?�?�(��`�{崱l�]����քu((Z�����y���:3�� �K����2f��;�HT�ݢ�k~�`Khl����έ�d�5����,K�525��Z��.K�]1Xo<=�&�t?��[�?�Rh(��ϝ��&��wJ��`��]�Y�V>Q�G��RJ���ٖd�P\�<y�O�'����M��-������\��@}�q�	�3()�����+��ئB�	��F��g�۪l�#Ǒ��Bl�09_S�UvJn??4�^��H��m��@�} �0~�N��ͻ��]�/"�<bW�Xe����Q.��ok-'���H��ѻ�9qfg�9h�9骜:�urx��h��5<o ᦹ|3����{��	_K���)c��כ7�U�7�[Ѣ?��3�&��~���\����X&i��T����9ݸ��T��p'�)�gx[�-�T���*��`g�-�������d|� ���҇�7q;U/C~���>@ģ������qG��9��V��U]���ncs�=)�Q�WZ�2�X�$��i��Z�A���>�Kw����%�1���'�|�R.P	����>�]�7�Tw�]��ݞ���n������r��T����<���S:!�4�~����rB,��� *<Pԩ�ϲ�S����G{��#����[�\5���)K��Z�y�q7�_����\�w��9�����V���Ԃ�y�a9AYy e}C�Xv�]�7�$�~�E���k�g�,񼶿�ܶ���¿XL��.N�qG��1�+5��+%�q�C�/��M��O^��_|P�ݢ]K�e,˭7���U4l]��I���5�߉Zf4���=d7
�v�bpw�0o�n4-Ő�7�
��Xl�_	��h�x�S��y��N)��^��R�5A�� ��M>W�)�:��%�+��"�����A��	X��e2x/|E������h�n,7��������_l��Ӹ�{Z��ٝ�y.M���$_�k�^6������~^Z�lOGk9�,(���^�V8��g-^��R?�K������vw�l���DTr��|�͘��k�M���߾�Rؼ޴�T ���K�M�M�>�b��W��ڷs~?��	,>�{FL��N[�ď���B���|��u5�: ���j�IWs��F�T����$|oY�?vM�7�l&�������6���kB�3A��D:��E�\bj��JD���M]B�Pϸ>�7U�5dv�q2�}/?r�,��87j>33j�hᖷ�Y��q����]��@�)0�. C����<����t;t���޽����uu�#3-�)��Lc����%�NX65���y��O��*���;�rB�)1^��k�h<E�dh2���K�IB��+5e��.O+]��Q����� ��nD|{A���?Ϫ�J"�'��G�������|R��T��|�
���$�{���$e�1
���X�SYl�~N���l��K��$�ŋ�*��[ș�W99
�<9�����9c��S�L�yL\V ���SՑ������hi`�oGҧŐWܑY|Y�[Z=�D�c�̷=��������9��u^�/�Zi3}���k��&	�ux���*�S��/�4�c�}�X�ɝ��|��f4�9~�'�\;����$�8>*IQ��H�&�z��|q�{�pC���ܴf�g��3	�o�Z&�!#���~|�O_W(u�yxk&H,�{c��ļ�k�M�/����љ_���[���^%?�t�)���|j)B�f=�l�qM鄠��sO��*A��������ѦS��MX�;G�k`$H�Pf��Y�;~��b��>�jl~�.��:���}��~�,5�mLy8"x�(��A���!��{*4�U��";��{��>�K��]y�k�a�oʀ�d�]���"�*:��#��F$^�C��+�jI��f ��u�_)d9�'��7dm<NY��f�z4�����kp˶pG�&$����˳���w-m�9WH�ϐY���yR6��(�rϊ�e��
��"^!qY�j�'iO�+=>B�/?f��-����̻���!����?5���N5v�>��0�tKV�W��fl��Z(��n��6K� ڮg��ml�yJ�paK ���KS/IC���{hz'��-[	��S|�R�f���9�z���ȅ�>:�,z	>+IjG=�Y���YH���>���߄8��������qJ�6������g�]oD����0�p�^mQ�<�zH�l�/�?l�x���P�Î��5���W�9��(#�*�D������)R�ԑ��H�V��Gy�!?ڷ��m2fu{���koh]�.ɗYI�Gu~sTc�]�n�������ܳ�	�;��k)����@/�F�;�JБ)�%��pj�k�s[�qn �d3-�i�n�G�J��7213y���Q���#Z@+jN2��bj�B:��IX&FZ(6����|�M�埭�����v�����A��}!���%l�޿�|N�_C�A��qy���#��5�WhV�qr�����"�C/����m��Ŀ8�|�Nm�ſ�������$�ș继$�C�ď�����v�3����P��#ߝ/ԇ�X��0Z*�ɕ-4߄��~��5���SK���.{jh9��c?�W�Q��>�A�*���_r�;�:�z�#��o<������S�C8�8�Q���]N+�m�?X�r^"pyH�E&�(䬎�/,���k�:VA�r���_a�2��i���N]�����6g�"���*�}�m�����*��$����Z~�����,��N �׸-۰������<~?��'"�٪�����7F�Tg�ߺ��h�d��r5�����r�-���S�+-��,��zB����l/�r	�[�#�vħ�&��]8����#�͊b��}y_��'lx��I�yG��?|��D�����>����&�����zs_8�����V�.͝�򽒴89���Y�-�f��E��MhFڻ�U��|�MO>)����s��H�Ƚ:\�M}�r��Xm3j����a�<"��%�%::�J䓠u���=��n!�f-m����ו[��Od@ׯ.��~��LmuV'��%��z� zH����DpѪ����B�(��
4�z]D�cߛOQs��<��#�Nn�q�P�����~��0)�֬����`�05��6�0]f�c��D�,��D岴�����u�u�?�5qo�H5f�w�SgV�&3e;Q�ٌ?���̔o���<���fz�g�搈���Q����>��%*��ѕqCQA�����N�m�r�ExD�=���<ex�M��r֘ͼ�^nO��2��`�o��������@��<U��&���v����0�7
k����1^��Ch���f���g]ؚΖ��9?����+��;��3�k>ʌZl���ȹ~\��HQ�߁��)������_�P��>��K9���R?��Yȝ���w�>�N�&b�"LC߻�^,�~2��=��h�ǟ��+��26Gl�n:��M�k�&H�
��>L�:�5~(vq��{iE�ûz$��	I�|~�4�{33R���[��[E���gf��>�f�^���k�ʹYM.����G?%o��<�`a��+�����oP�P���>�伢*p�-a=MH�5ٽ�z���@�IA�G�N�w��du?(8�����:	j1QŮ��g�
[�9�!%�'K�~��<���m��ȿ�����j������*�D�j&��Pߏ�"Ѣ[fK���\TU��17U%9�%�ػ�l���|m��n��F�C+p���yDw�,����s)���Mw^$�a�/#��7���O��� W{�M��7bq8�����o�����t��Y��k{��i��g!b��"(?7��k�m��1!�+�1�[tr��z
�n.��q3�o�=J�j��uǋ��0�Q�{Y��ᨪd�6qr]�;���/����{ϕw�>�	���Z�e�X}v�n�0h��	���M�	��`z	�9��]�ꕟ~^GrvEl��[{{V�o�L���J?��#>�8<{�0Ԅ�wo9N3J��йH�ћw� .���xE#hzdHH�ݪ�������jꊦ�f���=픤�A�]U�]�螰iȒ�����ެ�m�k�I�NZ�ʤ'x4<ڧ��x_�w���)W+-�$���I�˅��B|�����Q� Ғ +3��E��r8&tӶ3�����Rڡ�)?��s%�۹�,u��ׂ��ئ*#�����4<��L����gMfV����+{��R����%��R��Ǹ�Ko������g���CL$q���]Q�G-�'g�M��a��+��F��Ê�{թ�}��ܿ꠯	L�w�5����u��D���^a��5�敗[�%a�����$&����)�@w=�	��SpAȝ���P-����_I�3��w�Ei/5& ԅ�_��x5�B�\�E
�iߖ(��u��}�^������d�a�F` �q��I�~N��gf7h�%�����ȼ��=����J�~yڬd틏����S�.2����zorDN��N�d����v$껒~b��� l��9�M���I�gʋa���R��䰮-�3�^�O����{iqKӶ�3�!���{śZ�J#6�?4Q38�oE��7��O�0�#�"�6���$n��.}��(u�r�v�4�#�}]S_A�����������e~X�2�X�ǺK��=���^���G8�%�Et��ÏۘD��	�����~e��4�|�m2e�ծ�Z?d'�}�p���hz{��2�\��F�HӚ�%?V?mO���s�:�y(��~y����x:��3��gN4̖[⚽�蟱ۮ�ÿ�Y�8����9��+33:�yE�{\�� :JN��o���ãh�?�<�c`(�+�ߙ���X���]/���i?~��N��A�������[F��.��G���n4�>EG)&oS�T��{��xVh{���Jb��h;2���T�1.�@&ح$;z&�ؙn���M]�c�Wl���Y|��Rk��Y'��	ݾ����=Uw�^ׂ���*�A�J����2����Y���~���Y�O�~m��9{2�,�8���t������?	;>ޝv�=	s(�����]ے���#z�ȧuF%���]q��M�lj�hv�-��ݧKp�?�,��/��J������l �F���߽�����pЩ�a0�!ټ,."��A;��Skr$�<c�Z+��:�7���
��/NT͂Fga9�T\H\��ͯh��9о�M�Ѕ�Q��]��)|p����|ra����#�]9!��!�dQ�J$e/�����V~bGN?�6w���=�\:��Ug7!Z�����]!�7_�(�|�h���/�J?�PT!��ҏ�Н�^�	�w���=ꡪ�P���UE[��1�nތ��r�>����N�s���^�����%�R�&�]�Ba�-���Y���_M��|t�g-��I�̏�'�f� v0���l��Br��к��΃���]ov�hʐ�ùkR�v��>[���f�"Ύ�N�����L��+�	Y���s21o ��nX���o	{�~L����6h��I�1(<Ҡ� e�SCRS�ۑx��x`moʿ�+7un��&+�.��xCȬ3���f����+�k6����"5��7p�-�8�}H���1%�գDnZ�)5Q�	(��*�"��~V���S�u{���1�IeDZL&@���Al�F�ie�E1�����cݣ�n`R�/�g������;����L�!�mg��Z�8����$W*�@>��M�)���t�ʊ�DH-XeF�v�7��_�E�UTKXI��_�>�#�����
��@�f}9z��6�]�k�Q�|��	»u�;��K�m��p�I9v��m�zR𑫞qG3]}�nbv�d��qY��괯�Xh�����ࣻ���3���v�����t!w�ɝ{�5:��ˍ����ן�H?�m)r�d�_'��#�6�� ש�S��>***���1JRYIֵY:�1�	�Ν�]r��d�z#�:���N�$�Ɇ*ǡR�q<�N�͹ȍk	���Q�����/���{/7�9�N�!�{>,1���|�G�̃�����E%��]��zpXq�� �#>p3�݌�i�#���/=�ߩZ�9S����,��{�����|^�SH���3����3������T��6n�ߌ�м��� �*̓Ǩ��Ap)�����%/�g�h������i'c���_v)J��(%��L^]{AJ�ݮ�N����Y%ӿ�>�V��x7(��:���K=��4R�!�+�ͷ0F�q���$.�ܜ��c_�^b)�Q�F�Q��k�=��[���#'�;�#�H`U�/�<2N�9�ͳ��������g�����{�(����x_��Ŝv��B��浶FPr'�'���%�t�3�T������,�)�]�P�,��䅷�?5%yX��m巊�Qb��xb�]6cbX%ZɃ�&ݣ�ʚ�>���^�Hjː2w��^h�7 Q��oE9 x���3ڹ���u2�5:���A|,��!L��¦���7d˂���2D��qJ�s��7�fX����I-�؈��E9{^C��	�6+�ԪLW@=6yu�s	�:��.�Лrl�q��w��E�L]���vѾxQE������n�����r��腞Glo��Q�K���$�źe��MF����̏��hK����I���>��muZ�g	j���	���4�{[�w��޸0oJ���`0[y��)��h�^ȕe����M�{gS!�_E�Q����mO}yNL���8Б�C��92Ds���/��ʑp�4��O�I*r,��ڙ�Rc�U��傓K���%^�ȏSl��A�u������f��^��)�[�׼˔���{�ŧ}b}n�E|A�Q���G{�`��`m�E��K���R?O��ys��(��1D���{غ<���o^EX-�版�>�xkf�B� ���h1�8:�gq8e�M��ݦ��3-x×�X?7�0���^�@̗�G(�\)m1Z�M��"���D�����@��m���ƥ[>��y];�u⁩��l�
9�aD��g��8h������lc�ݶ>�ZmMR?+����7��^=J�=?%�������v�u;���V��xxw��D��N��T��gg������`@�r}{|�3z��6�t�kB����r씀!�Pձ�o�:�m)Pv�`����Ak�����_���$v\�[���ee�:�K����b���uZ�'��іQ����o;2�bi+ē��,9>��	�m���q���ס^	Pݕ��R%R�HK�y���45Kn훼jA~77�:3V�Hk�?��*hζ^c�7�G\�W�H�_��"��א#M$�;���`�?��Plȟ�o� h[R8�&��Zl��X�E�����&޲�-L��[�pؼ���_憢��F�����:M$���q~��E�������������%&+_�?�=ݸ��j������@`T�x�B ���K������+}GXv�-w%����܁L-�����G�����!��ε[1W>o�^3�--#f2@4��tp�����2�f7qy��oQ�h�m��叝b
�� dN��F�Q
�Ϋ����,[�y�ہhF�Y�tt�y4����׊���5��oodi�_����wU�����O�o��M�o�����V�#�6\E��<�=���5!��,��.'�_�ۙ�W/&M�0��ד���U�qo|��xr|(
��쾃���]��9N�l��K�n>SU�1Z<1ߐ��K�J��U #7v�|��""���捾����d:Å�QJ��[�#m��j�Oe���.k{.��dΟ/�ڄ]O&�>��!B��n�GD�s*�gz���Jw�AM='N�?H˛P\�s�u�<���
���~T*���&�#�o���������_�#��S[�:o�U�A㓨<7l�AJ���/%��?�lrz���\ߎ�os��#��.�cz�:��!�ɷ�H�Th�V?L[:pF蕍 ���4Q���д���l���؟X�D�2^U�NF�����St�7��~z?y7q�����N��u�E�6u�t;��(�������g�&����XDws�A߀W����,�K+r�S�*z���(d�w�����<8��VUc꺄�ל��C�䀖�l7/��j
�xְfA�d3c	�>�)>�y��^��/Dz����MȭR�����a�'�BG���=_J�!�S�grZ	���<�0��x#;�IPV��H&[���nO4k=�	 �m�W����N {�g�N��(p���M�\�C-����t� Q����%N_J0N�S)l#�U�f�d�2�R���ҁ��;oH�z��7����ʃD��B�ฌr)��]�+t�X]X�Aw�������>��'��������^3��0��G���		�����X�9A�rԵ��یi�}�l\��jU��Y�^^����ne�$�0��y󆜾�ǆn7�,l���=�����4lty����S����*=m�"C�,�� ^�0l�h��U��G��$�OQ��6���	ؙܼaJn�z�$�A�����2��eɤ���L\�0�˺A�v���BV���<�C/0kiÒZ�H8D�K�5�p������������|�/#Ò�}{�'�3��i�C2V݇���q�L-����qN�j\g�r����H=ч|<f��1C�$k�'Il���0nW9�n�rx�./,^V��7Қ�֯���d8������O����{W�x/�*�Ȥ���a:-Q�Ƀ{OS����<�tݣ��/�i%���,+y��������⧴d�g7�{FTɗ���ޚ*�&�L�af�;�J��QJ�:�;��賉��3zX��-��e��>h����LQ��7(�S����J~���Se�H������ �>���?~���eԲuf�-���Y��!}� 5*��D���88�+��ܵ�Gkϗ�E���tI�5K���JKun�'%�����杢C{JMZ��Ս��jr����W�6wqf�n��r�5#�gT�r��.:�/�J*�ߩ����?�j�;�����V��զ��i�}�M�4��ȭ5f��͟��ICY,��2�S�g�^l��oؗ?ٍ)��ltSc���wV6��D���_��u���Z�|��|�t?�i���i�Ǌ�#�+���\���"��ݡ諯����-F+�-L������"��;��%�7�@C/�2�Qc��c�h����{���V�D2ٮADe��Ϙ��Q���;� uC��+�$���;�sw��4Z��VYwo�Ú�b~4d?��ǘ��޶#zM�W�|2�3��{�`��ߧ�tY�\��+���+؃��a�|3����YJu_��@�GG��6�����@�撍:�Xj1�_��.������E����A�
�ao{�`�M�\��G��Ӟ_�pn����k�WY�هV��ڑz��\�Y�y�~|��Y�Uˮ��E��a�}��a��J���_|��1A�Ξ�ށ-�8¡��ݑk�>�ׄ7��@��5Q�wY�����6�,'��!����>����״�z�v�[�&��JR꾏�*���Z�8k4�TUXh�b^|�HI�ෝ�����F��ɳ#�\�=uγ���x��(�%�5O�B��(�Ѝi����3���F=
��0��,K�Y���]�����A�����I�&�j�G@�b�(��5�p������6��K���b���� �͘�x��_f�Ӻ`�}�.q�'WO֮�D uk������s�.��*�)����nS"��lj��Y�L֝��q��u�N�Cv7>v��yAk���~�leV������Du�n�YPY<,��q"���-�^���m�=���<ɇ��
����d���៱*%��&��(�&]� :؛�M�??,_c�P��kG@�ق����x �7}a�!<F��Sezp�o��0�uW��Na1f�8ŭ�l�E���"J.�2�;0� ���	�M��N}k�Y���ɦ8J�Ȧ�F,4,��F���([-.K!�ße�.�`la�G��hW��'�)�&��&«PSp7$�����gc�M<p�U^|,�&+	Sa}��i��P4�~C�4��
���u�5���=w(���yT�j�wg�-��]_�Vi`��䳏���
"~�9K�E�#�������߶�7��q�f^A���Qv.�Sj�Go.�ng�V%܆��Q`+��$�誌v�B��:'Զ���d�I�.��T�;\�q��T�{$�e�5}�r)U�����0|��#8��:Kg�/c�e���V�.IF�i��7)G�r�����Ƶ�����D�"ŭ�^K����>e��5�'��W�)����>k�5m�Z��_��p�1{21�gpx��=O�{��WN�t����փ�h��>�F;�ŷ���˺໿��ؠe��=zޠ�}h]��w�
�� ���@�o�_�00�2�0z�К��x�>I߃V�̗�1��@��u|Y���h�xi��G�4�c���c7�yū��c���n��K�n�E4/�~�|ȕ������kT�Q�{H�)S����/ �.��6�p�G[��R�
�C��4#��I��v�C�iu��_����͚]�{��UY�!�?����'#0����?u��r���ic���LͰ���n�y�2�o����v�e��n4���u�]pM�Fҷ���������p�*pf6ҥޝ�iw<�_�%|��+"�����1�'_+��t¥'�bol��K�UI�p�7�C7��Q���}{�?���:/��j,��lP[��.͌�m��:F�_�CluS����/��ZSZ���~\^�Ɣ��b;
e��*�P��
;`6'բ��?-�s#���KBf>`��u��?�����&��1�-/ߑ���&]�<k�8�7�S�z�$6���y�,}��~\�ɡȄ��%�G�� �'d��?i��}�C�^�q���H��)���9u�k�����B8\��pX������j^R����a���1�Ƿ!I4`�iY��U�������"^	u���<��w�6M{^jT7��tC��L�����k?O���1p)���"%À�D��8C��o`kv��*�t��H�
󙃶*o��Od�B{b�^H�k�M�c :>��zЦ^��hv��$0��s_��u�rX�L��+@2QXa�[}��
�u:=�n*�l�-��6�P���w����]��V֒��e�Y���M8����C.��[zR��"�_���[����� �����|d���.����H�bZ���}*���bI�Z�����Um��.1=y>}J<v�=��a6��V&_��d�s2
C3ݕ��#���y�SG"o�2l>͎w�՞_����������MU˼&����4C$)�ڢ����v�M�i]eP�������"*~��ܤ��8�����:IH�x�O�6�)���U�k��)���U}��I��'�#캪��m���+�o���ľ�LGl��-l����[ay�z�;�&��ʽ��ؠ�S�^���-4.��\�`�Xҍ����	��Jy�"�SZ�IԱ�xK�H��������K���W!Z��6:LQ�6)ST�(�طXne��֋���i* �	����T�;��ʪM����0
�π$ZG ��;7�kb��E����F��ژ�MN��K�K�p9�U)�Ŷ���bjAX?��8N>��X�]�~]��V)�`�O,1�H��ʷ��~�o:f֦wK4&��f\��Kj?�R4�E����!��U;+~�W�l����vy� ����FmϞ����;�;7�АRV V�2'�xtc�Z�Q6itGU��$�s�#��X��u��1�oe�}��
�X��������{�c;�tދ�<1<�؀U����<�ˀ3�q��Jצ��ےaY>�q�Ȅ��7�x,Z��T�=0���2�[��� rvYw;�8t�ܧv;�٣�k�����}J�z�,콋��a���("8�I�,�B�`����w>���5���n�o�֜^���@[�,�uZ������ܭ�	t�<=���7�Mj"�y��������������2�'�'�"��2���ʆ㴓���{y��Q��2b�aL؀��Y�w�	'ܖ��Җ��$���Ůͥ�����j؏�{�i#w��A�^?�{ܠ����C(�O��b������:��q>�T[,���`Һ����Rʵ�S.+M�;��KwQ�����ݱ�oG��a��y�.)�����H����m��\r7�c����D�H����N�����UnTK�5,�xE��;���2ҟ ������G���Rg�U�<+o5;�k/6q��:ݴ��#��r���b�$���JP0���.�T��e�a�▐Nr(��D�_H %Y,�aIMw��'�v�8�r�z���/0蔰7,}m\75U���2��TЂ/��9���P�5ڌ�����l�����=����jy��'h���;]ؔ�� �z$�j�����د��t�<ڢ����V�׽ܹi+�������y�%��
�`L�G��9<��@�zݠ -|~�JPms�|�^kR2#����]$������S[��t?=u������k�M�+o��^
�^}r��9��$|:��@۷���q�_A���2W��sik��0��l=(��&n| �_29>; ��O�/C�/5;m=�62Us� �y����7sDv5?`�9[op-[jn�S7������w̸-/H3R6����j�d{�p�(��6�G� R}f!F���q��������Ֆ����]ǳ��?����6�bMFMT+��Jy8��;�L���������D��jRE�q�	+c%0+�DBa)e�f�o��*��3����j}Rb;e�'�l�~���Ȁ��|W�
ya����S"�cR��I�"��ݲdW����<��� ���Uc�&�d����Z��)f
���8�dٛ��@�2=ʍ;S�����#��,��R||��.�=�����a9�å� �����yJ��~]Yx�Φ]�����k&�Z��&7H,�{���욎��70� f]��EL��/�DZvM��E�K�k�T�;lD�S}�p����!�cvJ��ݮ�H4� ���3�L�J{$\R~��5����_g�>$��`������`��Mٸ������	j"� o��۝��mf�e��L �.�C�g�ȗ<��2�F�ⴂ�y��d�ǲ'��\Bí:�V�,� �8	�Z;���q��t�z��L4�ʈ۸����\e:ܨ�W��++�Z�0!zC���|X���	��`o޹w��v�K�X}m��Y�q�V�;�ذ���f����[�G��[��N!��9x��ES@��)��T��]�� ��˙+g?˔�8�rx�9�G��2�}3k/�%�L������Gh��5�l����������I�e�$C�B�v��穒�FU��?l=������;�/?�o�:�b��@��"�� ���!�%S�-m��x�΅�k�kf��Y�]��r��*���T�Phc��7�5~��Q��w�;��������Q?�Ll���u#Rv��}u_<��w�"�}�Z�)r^&�y�xlЎ�<k��MA�^��w�S?Ψ<z3q_�{�-�ʟ��19��קK�T7������/����$��9l�~�'2M��m�A��������fW�r2�j��T���A�F�L�%$D%&w��X/ٰ�.6&"ʖ�ꢽa�l�#/F{�?<�v�H���a�m�kC�e�����'Rk�THu��|���
un�U����畓�(�
�O@�i�c�._$�d�Z�;bxzz,����"iQ�A$Z���0ȺOY�nÝn1)	oȐ�g2j%:�
�<�̈́����z��V���2b��;���7��^X��#�gJ2p�nɅ'+��tn������#��� �>�cf#M$���-J'7t��9fAO���ߴ��,4
��z�)t��`	���S#*l�&�+9;H{N���N�>b@��.;�q,��F�r�)�o��߯���.��2&��^�C%���k<�s����k�n�!�̲�>��H�e ���N�B�VAt�{���s�/d���I��d3&�ƀbC+��~]��Զ ��T*��~���*���²7��Q~7��0���*"2�<�4��L�/�z'`�x���^;>�53Gsd��65Ǽo�_R�^��p=�J�栺w����E�9\A	M'*����"��6�o�q|���1�"h
j��� 	%M��-ux|�SļS�Ǆ�o�RFJMd7����h�������*� !"!�Q*�#D�;F��"!H�tw�)��`c4��F��?���꾹o�s��s��ܧ�8NH�u�+^�U8Ї���ޞ�x>� ��u��}��@6��S��]A|ו�Ƭu��e�\Q����%�M�Խ�5w��b����/znY��&�
�����÷����d�C*&!6�� ����Y�GL��\&E���s� I�g��Aܾ���=�_�=�F�z����J"��ȗn���0\3s���ٔ����T[[�bt)���%�\��z�P���'�Z�����~�.ͱUu�8]q?Q�j�-9J�A�.C������s�	h�w����7���o�	Yّ�+�eOu���p,%q\܄8������Ǝ	Mh�o���l��0�q����i�|�&O��].KUv�A�f�r.��l�j�����wR��/n���1��0dn����)4M��\a���g��q�M��j�/��,N�oB���Ux_�@۶Ok��ټ�֋�Y�+*2:0�2�T�K�/2�O�B�dT�ֿ���
H�LP�7�rs#�-�{b��#�(�e���YVÚ��#��"�y�fw�ƾe�P�Js�@k�e�NO����~�{��g��3�l�l��p��Lѓ8�v�e$��)��!�N���K�˹a��E��
��|R���u�T�?�.�6bȄ�O��mS夂S
����dr<4��TC���������2�v��'��-������o�g�N	�fԿvl�wJ%0�]����cG��Yw���M��r=�v�ou��qo���9�����{}۬���ݛ��ʤМ���C����vڂ�KN5��Ȇ%�+���/�}�3���װj�"72ec]��r�織�~�ԉD�ȓ�~�P2*;qc�� �5���(ě�++a�!���8~5K����-�&m�AB9��T�Y���Ag���D���?�p�����T%�����jl7��v<��z�ݱt���|XC冚./S�t�Rdn�
��]Qj��	�]z���*���k�Kɤ��Ȟ���Q淦f򨽮LB�{_C�$���讽}�uGA�����絮���O�|��-��9�x��Ũ&������b[�Ƅ�cO %I�W���|��r��C��<f?�b�����T��tq^�h��N�m�} ����%K8D�E�agl��be9aK�K��#�2;sՄ��X1����-f�BŒ9��u��������-�V��4�Z07y$d7��r��57`{� !�r�Q`�L:�n?S�����#�㗇=����MɦI���Ղ�iz�_��!Ogf��[������rO\������L��um/�om���2�^,̷��U�>�~yP�Z��Kd�[�WB�Ǭ�)��q�K��|��aZ�9*�r�������_�+�1�	�{ꔡ�D�I�"��K����Y5��B�!KR<Gz���l$["	�f^�?�+�e{��q�ԒH��h���շ���C�/r�VA�=�c�*�;E�"K!�U:T�R,]��l���$�d��7G���n\��8s(�о��4`t��'�;�%[�ې����-�hhE���A	=``��U���u;�h�Ϊ�VYt�x�z�]#o�5�e�	��*�͸<R˃��'�U[~��憼��ZRB憖��6��΀�F��BD_��I����r��
��G��%�e�\Fl[믇��I�Y�7��j�uTj��v��?I�6DN�	��O�,� ��$��_�@L����';x���n�6(���r�;B�@�s��mƻ�YI�O��s{M�..��讻)"UP��s��Q�A�ee(����Q�d7��QLa˥��j�&	�:N˦��Ч]���-~���!��g\"��\��lZ���G0�ӟ)��>��e?�=	��oo�90�)t�Cַa��W� miK�R�U�5s�w.*Mi�E�Aؼ����J�P�1�	��YH3��v�F$Y�<��#;|٣Q��u�]�Pȗc���-`jx��D�f��Y��isibg\c�ڙ��T���7��m>>�XC��,Ż�z�`Ɲ?`��"?Ǻⰿ��_w�<4=%m�`t-=�?�}�׹���g��r�5D�^���7?l]���������J�-�I�8Q���N��ɷ(yO&��O$m�U&t~H���[��>�Oξ����-1I��E�g�L*�<�q���=S1�hY�ίv�*pe=�-$�����7����U�	w6s�������p�j�+<3�(�]���ڗ<(�3�|�o]���r�YA�%���I;�>=~J0=�C�u��q���_��O�I�)��TM�
+Զ�3o��x�P����hΓA�G7�BFD��
¶�@|����/����T����wc�c���֋7Ĩ��Xqq#�[��o�I܄�_k�l�&��~�+)��+e��Y���߶��k��n$�=Ǟ�y�q��)��lM���	��Ϟ��2<?D������O��NzY�H,�`�xڃ�/�]C�z즎� >��>|�GM��AǷ�\5"̋�L�a�r�GzfR]�a���"T��gk�pƙ:�m�={"{�_��6wk�^?�/,� �jL����]��%�+�n%�<�pf]ᐍkE"��O��*r|-k�Jڰd1�x	�l���]�y�H0F�'8��9�z�oh�oR���j�ƺ��B8:Էt�g+hj�5��"5<��Zd�81�;j.��!���V���d�E��\���DG-7�Y�2㻦�2�
8G�b�ٽ�߳�ctS{��Rk���R���j�z�u��gi��^�A9s� �<��t������z�ԡ>�ͷ�/}p�
mx<b��3�8 ���p���B��d\n�4J8C��B��&a��N/�39v&h>�g��=����V�cl�����5+�m��s��׷g$�Q��K~D$	�n �r�{<�	Pf^k-(ݻ�T:�*�r�����\6o�4W5��E�Hl����~`���)ʹS��t)aK�was�#ۯ���w���8�E����;�j�wA'�e�&��$|�V� C�Ki��e̒f,_;����z֦��@��)�@�����8�1(�ݾ�npʍ�S>|�?���}�o�����M�:�ؘ��ҡ��r���y���2�Z��\v�=�^Q�
������8?]��O��)�����H�Iz��ա8*6���'C[�;e_;ds<���1<��IO�t��y�0J[0Z�}��~Lc�S�{���\��9�b���E�[�^�η5K�q��]�D�b��;g�\����sbbj-{�8�ӳ�'��� �uK�}��F��*�%��c8�k�/P�1v"�I;����E`��!R��%�Ƕ�ّ� �5��b�Ik\$;��Ġ�S�����Ҷ�� ��E��;�_Z��w���?���[�����-�»���<�nr�z[ћ��2�}޿b��m��n��Z���qn���8/9
��y��z�W��RQ{��S����o��R��7��A�5n�Z�l7��rB��R��x��\h�c,���y8&U���B,�|��j�#�\a�u���9�����6�>3����_R�Ef���%u�&��1�.L�'n,�l���P���5�Kkݒ3�#_KC�u}"��=p/k5c�!�?�*Mv����Vܿ<�猕c�: J�KP�WvSKY̡��9-�ҟ��_�����7o�Z
�a��\;u=�a���|U^jH0�ኊ�f��9(|a��/c�k�<�n��3�R�,�.���w{Wv0c����P�k������ת��Q�.���`{�W6I����, �	����t�/tg�	����Ðz�vA2}h�K�Ԥ�(�@6�R��*�^:���{z���	�R����6juX�?[�P1��"����~�^I4w��!��rd�����j�a�F�Fu�a�Z��|��
���L�R�.�]Oux�_���������I��^�]+�?�����|��lb%V[@��i��5-���l���9�.��$�0���~ܣ����I�h���t�y���{_z�@H�b7��P.w�p+���zI�ܤd�;�S~v�ǵ}�[�g�.�t�ׇR2{C��v�·!��m�����l�vf�?��"z�m͙�'��/|�fE�Hx�vC3���p~�`!���5$�-�֫���Hl��y��A��%���eg��T��)�O�.��`lS?Uũ,DMT8�*�ٔ�6�����і"��
.)�?��1�����H�!���s���Ӣfz������r����X�1	i���ՆS�SCU�~��q:������T�+�Mư��d�y���(�Z��!߾�T4�����N-�v�1�t���OdRq �R/�������ˑ,�_é�@�cְ��q�o��ڪ���r�/��V��%���8S���g�������D��h�1�uP�����{�﫯[Bf��.�[�jj_5{&]ߎx�=T����*[�Pe����L�؍eH);5+��0ϲdr���B@�����*ҁ�HO���<(�`WP�o�����&��JS-:ν����*��G�1*�o����o��Y_j�n$�(T�h
�Δ�}8�Rj��
Z�mHD��5; �2�k�0�%��nD����j±�H��jw5�;c��R�2� �B7�`c@��X
�5���Q��V�$�LI-�zOi�y$Ԭ�����'����1�^}W����˴<���T�O�����܍�ۊO�� S+\n�3H�i�釞�qRv��é������{/���=]����m����,��ޭ��7�[��3���!~3Nl��`�j��
:��A�H�?�ژ��̰�9�j����xq>�W��|�p��]�<�Z���g�Gl*:��3�U�?�`�q����$y�]a����yB#$:5�3D)Qg����rLט}���5�=)�����r�� ��Z�',����a��d��d�F��y�k��3V� �:\��������w���adl�/�}��� 8�:���JbY1<"v,��~��xp0-�{�y\'�JA� "5,��F!�迺�1=i�۳Az���@#D!1��]�#�b;�����g����#+1ݯ3�q�(WCbu���+��o_.k�[���ʂ��Yg~���U9j]'�魙]H\�o�J��~	�yd�����8.^��/̳y�y`B���2�ơpu�g�_��s{�����ȹ*Ğ�N�GcImg*i6��		�)a��H9����󀡖���b��20l7�Z���&��p#:�.�Z���3k�&��T�{O���.�N�2`񚯆���%ݘ����י{y���.�!1]R2�����]*Ҏ��]�y����u�G�O|8�S�a������I���,vֶ>w梏ۓS�����s=d�:ku���ۑ���x�(��-9�%���o�/q��0ȯC���$���
��U�r/�N#��*Op���	"4���95b�<��w��&i��d�ɨ�Im��<ҽ�Q\>(�t�.����A8�%š���Ecm;"|}}lb���>��^���:���}EQJ�ԗ!�`H�a㑻�B֕ʱ�%����<}�M���<q`I�g�yl�rxߖ�#}0�s��$�I1��E�������a�T��0�ttB�|*U_�Va��������Ql4��n@�G����ՈNk\���� �� G�xr󰳂�� ���~qj����>�i�j5��k���Hq�sG�#��+����케�[�5��'�}����ǯx.۶D^�Ll*�֬��؇	�н��ʎe����F��w㹛~4�^�Was��$��)h�4<W���Or�%�n�N����*�]�41�� �GZP��/�8�"�5��8�{��["��O��ȡ@�]a�{�F��(���w1'�8���=i����������'.�pķ�"� փ��B j��+�@e�ү���(9;�����t&}g���?�~���o�{@d����x�w�Qqӕ�W��5�p��?��;y���T�"�"~���^����q�����{b�%�b��!-�3�Uxx��Bϖ�1-�<��6<T*�J����
�J:U޴&=�ҷ��|�����e'X���z)aPy�5w���i�2�Y	��X�"Hzɐ���C���u�sB�	X����s|��B�$o����od�$oK���RF�O�ei�	'�F�|"����-C[�������q�؜;��}��i�!=K�W�M�#������к�Piy�-��8�t��N	M�}$�k}����!Ԓ���C�S5nU����_+֚�{�=��7�|y]�zݼ�l��م\�,�\D��-��0)z���_лo��T���A]���z�};��l��ܝ��ő
jl6Jݢs��( nF��ط��R��o�${!m�n�v�S&���5��(��/�U� ���v�Y��YE���ks\�c�7ǻ���:�)G ���� �����ާ��8�Y�;\�T�3�B���t��̏��ȱWt��Đ�Y�4���ݎ��L��� *_���N�:b����dܗb���G\�9��� �v6u���'4�Wd�Ē��.�)��čzݎ,��Y<e���(�����PP_�is2�%�J��5g��]���~�� ��;Ĕ#F����U���f��^�����w%2�����ۿ�&��2��
����0<�����!|w����)�{�}(�|�����B�q�3h�=.���l��b���4�p����R�0��?�f�8͵V�$)X���q�_�es�)L'��>�&b��Ɵ�n��o�o-*PRi�5u+�y���>���q���JsοBe����v�u�#��R�7�d�y%o>��^o������`���L뵺�c�T)�%��aR$?Er� �G!W9�`n�"�+.y޵S��)�XW�ӌ�z>hR�������b"A�G+E�$�agxK�bIf��ΐ+d�*%rW��ON�דx�x�	��%��
oW�O��}�T��&��DfxK|���G�~O7�bE8�k�Z��g�i�����Y#��k�}����Ǆ���+sl�F7�����}�ũ�hНD�E(ut飹�<�:�5;�&Sx���=�U�(MԁGE~L��h=p\��+j �kZ����/��8_��f�%�����j�}�H�c���re=o4��&}b��,���bJ��JX�0���~�g2y�*Rc��<9�e*�T���Nñ���w�Ȩ�l�M}hE�!=��c�Z�5����Ժ���Ƙ�,�77C�����	ۀ�ˬ�w��eu�Z�r�5/m��E}��ݠ���n �����p���I(u��'����w[���
�d�ڌʞ�kl�P�3�pZ���N�<:8��!4�zy9r�����;򼆠��PM4���3�|��z��֜�\0��۝j�,�֧���N�Z�=~����
���(�E0��;�[ɳΨ%�)����[���z�8���A͎`P��Z5���R��0 Ҋ�o�G5�G2?v4,�(��i�?���BLm�|/:U�pA��X�㟐ʰ�Y������R��!b�%iS����m?��Yi �-�v)�`���[�ez���QY;֪��n�@W���P�Ox=�|(�jF�"Z��`��^ ���FwKq��/`�W�Y��*��ʵ�|TVgt�4���$+S�@�w¹�Vٱ�+t�i�H�>��yģR��N����0��3K�!�yrբ!u�r�<�~R��x�E�-^��U��3���W��*a������m
���
��p/b"ƞ��K*��Ec�P?�iΝz��U�+�ZA~qd%�'����ң��S�n�Ƥ֥�q��(�?�T���Ѻ�7�E�ѹ��6���F��F��|���V6��!	&r]��zsKa��T�v)T����v�yĐL~��\�z/�l*ۭ�. 	"�����_�Q��sޏ��&y��1w���)U�����{́G��y&���	{T�k!�rKHB��UO���}h/�Π�~�[	R�(���pX;�X���o�]��QJ��s�($@���,mR-׊�c�CKv0�<����ا���n~۠�c\>�j_�KE�s��Q������bO��7\,e�(��)�
H��]��U�7;[3��?#l���I��&R#U�P�6�}d�~��C�dξ�횥��2v���rBY㉍���/ޚ����a{T������X��Z-�F�F���D�������ZT��u�@�Q�������u�K�a8$֚ݟ?\q����T;�G�옄(k);�8�L�H�v)c˞<`��i<�%��|�sЎ����mV[_�Rс�T�A�6�4��$��wKZ���Vu�4'yK���ɦ��i�5�����on�U�{ͩ��u�[���K�
U'�J�I�@S��|,�8��	��E�����E������j6w6�T�� Og\ߵ�_��ߎ�G�|������e�-����	ѿ���N��!5�P�9<���F�F�Z�Wic���H��-A�%�t(��uI%��H���n#�t���U����.�|�8��4-�����:~3�K2��Λ�����߁V�����c*"~�r��&F�y`B��'�x�7ek�	�e�:���̘��@���˱�)�i�HK���[>����ڏ�X�V �p����z(h-�IA���H����`��V�bG�/�^L��ٷ�h����H�.���E?E�F�.����B�
p��	$���¼��0�gd�y��Y���/��W���+O�z�	��ΡR#l9VcDq1'��^(�6��D���~w�)r�m\۲3�j)��H�}�s��헝H]0����oL�:/��B�J���3�1���q{��YGv�f�p>��n���+'MD6��"� 1��r�0���Ϗ��95!�~��6	Ӑ _ô~�rļ|���I�/k_wH�L�5Nqz޷�6Н�k�p���:9�\�_�Yx�_IlΔ�[2 qӈ�A�,
~��iNÏ���*M<���nb�}�`�?�_�8
/0q���M|6s����ٓ9ʫM*:w�^Qm��)_LW�nL������iTt��L��F$_�j_��.uK-��g���}I�,��I��t���f�� ;|�W}�cƜ;�U�u�͖|�t���w��CD���G��z���L�"���	��B�XݷS������ε��F5�H�A�փ�9r8Ϗ����;���2>峃���hǦoЮ��g�"�1us�$�>�M��Z���od⮖��B�k�d��˵V��%�n�|��[�&F׸&Ȳ���h�1D4hM�By��E$\+M8nЯ��ް$#���'n))܎s*C�u ��raΦ�	�C1C��fF5�ʒ��:���=�[����G�:���u�(��qz��S��r��bs�D���V5�Q�.dvB����������R#�1dj��hr��������ɱPZ~�GN==o�,�R��^����y�T�(� �z:���~}sx\'�Y�	�l��!�yI�&!��/������3iM�&W{BOG���1]�dԗ�Y�y٬a%?����/���*�{�7�$vn���o~&�쉉A�`��o��8D����R=�������Tߺ����O���&K?����bݿ7�:W��`|������|����"ǳ��}��i�z�t���a����,j��z�h�R�M[$��_�/\�Ot���\��u1�H:��}�6�ZNؘ���g����W� �s���tb�xNd9;�=�������:���ѱ`7�5v�p���q�6H�ܨ���,ahɇ���1hə�H�"i>��O�Ha�F��IB�������1~(9����[�t9u�Z�ׂ��.AX���4M�Խ}�E�p��	B�%?^�� L�����Eu��;���쀋=ֿ8wp鈨�e�^��O�0��ϝr\��F���A��"�{��/�,�n���ˀ)��RU�7}�Ug��.Ó�����>���~���O�:�݀`��.7^k��p��@}��`�/Y�Y��2�>�������ɢ7���$���c	�Z�	��V���<M�>@E�*du-KM`k���I-[�c��*�3s���)�ܴ���y.��,S5��cf�9^f%@��DnB���O��/)(9΁B��8�[nag�ԧ��?F�$��V�K�9F�sO3R*�����X�%��<��ء�U~�`rdʒ 9��B��E��bf�}:Ż`�P\�+�����Z>h�.e�j�r�f�_�!���x>yW/b�2��S��KW��4`D�^�!*$Й�-�SI�#��`=��������k}KJq����	��O�x�P35�~�kR��)�+��|{��3V�l;<�^E� fH$r[Z$*+�w��=�+�ʀ��r��js�%KYU}
f�Yo���p;�F��&~ZmK �Ҁ����@����6�jP���0B�Oc�R0e�r��v��;5ydL���.�o������=��Z��A5�+G�Rd�V�NQ�$8P9W레I����c];�i��j����C�~��
Xo"�SP� )�
:l\��� ��D�5�Cj�V�6C�s�q�z��4N"q��z[	��v|̬�Sv�wi����
��>$U,%�jݱ!"d�$�5���#D$�2w?;dw����Y��_����|�#�a=_�x�
ɖ��IO�RZ�8~���Η6um�W ��R�y����˯N����a.�W�{��wrOV>ʬ����$H���9�}�)Gaq�"���"��C�e�m�8{�s���7�ʽ[��G���e���8�v��S|�Yl����a�z��*g�Wʜ���H�m�a�7y��ښ��ɘ�F=iy>�/s{��t�0<�r�>W��#�:��ss���A��%`q|�'�{���ml^�&ь8~52�ُ�ϣ����p�x�Ez(ϼ���ۉM�Wz�*�L��? �ٝ�=��j?_ّ�����]q��ݽ�I����/l�;io��V#�N��I�)}�a��T<�'�d��b�&Cj��|ᔜv��)��D�Z���P)d2��yZx������g������|�^����A�G��{���ƽt��W9���_P�t����iȜ;�`GB�'Ks��Yèo�vk�(餞z�s�k��/'��{������4nIv�l�BW�)~<�fN9<�XVk[��7�C�����1Z�ߟ?�7������&� E�����x2�wb3vP�@�lxʨt���T���?�4��k����⪙�^l�nLi�a�%���
'1�jhѺS�x�����p� ���xlx߀FO�����U�-�6	�W������GDйwV�y�Lz�c��`��P�U���洁�bBYdP�7�X>�v�ᱳ!>�Jn�S��;	���
5?q���0�w`wg�2� �3	��z<u�6^��x%��iYܘlIp/.%$V��Ф]�i�ُހ8��n=��V��n���ń�r�
�~m#�A*�nA��\Ʊ}<|?���@c�h�
:�ʹ(���w���K>��:�̊��X�=I� n�u����	Ah��[U����M�;�vJ�N��[~��FV��N.&���G5�[6T3�wxd��N`7%��"��z�0�9U�#�߰Cu�i�w�>nS�Tz�C���"�`���3�h�jR�{�$�D͵���>��f�lM}�Q�p���1��Pc��F��|�-r�*�Hw��3����dϏ��<��vJ=4(v�dw��OBf���x��fE�Xߺx�1wB0�9 LZ�$;��Z���C6��q��~�dy��X@OTJ���������]�D���㧻�5H�0#Ο���1}`�Խ7J�E�0h#"ud��<ƚU�l�5�]뎦&B���m�7	�l�La�&�����e1NJV�S�!=m]~�Ώ�m��?�]���~�)�Rs����i��jr87k1$����Bf3�eYp���P���������vfJb��N�C����g�:ؕX7$�u�����J�� @�?�·#�M=:#{DҸ��M��|O�r���Ҕ&2���?�Uk߈����'p�Ka5TV9ސ&5w��\o�-��)�i�����߆���;e?̖�I�Ԅ��@��_�=j+��l�O��dC�*f�k��ȟ[�{�2�r�P. �b^������d�Z�0�Nm>��Kd�'uZ�i<�B"ҢU:��7�"SV���}�=vY�����vE��ZŚ�P2Z ��	6F*\�N9�ӗ� Y���lOs�{9/ien��2����6�������q:U�0�������T<؟i)h��Vz����yT��g��D)��A�i��ךr�m(C͸';uC1���d�2z�v0v�8�䒯]J(A�)��L�@�7Ц���#=Ӆ�h)�+a§�O�T&���z�vFCJZ$Q��Һ��ح��	"�����u�'��[̿��S���r8����^��B�4�M��*���R��"S�G\�d�0WH:}��x�-�;�x�m�}����܏�\1deo������%�X�uݺ��	v�_I�B����-��.pk�81-�ߕ�rL-#5dqՒ�I����GS�x��l�x�������Fj�el���O��Fr�!{�QَV�rӾ���AVv���p	`]��@�Y5�I�Lk����c�
;Hz�ô�n�K�MB2`}�h��s�lC�@zq�08vE��5��F�d��}E�4`ϷϽ�}f�N,��w�>��7}?�*R����Ua�(�\
l�pj�Q<�����瘲��$��Mr���3ޢ���A�;��"�����|n�-e��R��]#}M�h�	x/���/�U�Ǹ<<�E	}j��TЫ��@F��'m� u	[�yF�H�k��"�/g?��4�U������'��U̱�N�:s�"���e �r��w��=�A:��PY�F�f4�C�H���?��C�N��oĳ��c<�>�ɶ�Ea��<�]~l�m�l��Bl|B����7��~���ҕ&����Yz����H��j�����hd����(~$�a�(H��}�8���H^�����wD�?��5��>����ҭ�v���ܐG����9�;>�i5%�9�gځı�QJ4��)J
Ri	�ir���S��3y��q|�$ث�ذ������w�9J���[��T�a��y�W$Z[;#�Ux[,@�PC��?�W�!�g,��9쉙S���%S8Y�M
&�pv��,����A6W�A1�V{}�1�C���s�YhQ�(c�#�R9
�pD?'���w1A�G��ai
��3�v����s�zj� �O�Ų���Q��j�Đ���H,��T�s����꘾�SV��n���:��SK�[-�_�R����2���σ�rs+����������d=Vq0a_@;���̙��#Y�i�ɯ�>5�hT��[ދJ�E��9�>P\��S��aꭱf��^�wG�@D	�� pl��AζY�����--�Q���iS��8�@�s"��G^�3�Q���H�ani��
���3�4��N6M�ћ,6�5j���v�緂��{7�W��4�~�2ع��8z���I� [��I)�4�!H�L�.Cax8��arW�՞�ǵ���R�L�l������^k�xտ(X�~�����9*�{��'�L8�urS�J5���#�$,#j�C��M�Ss{9ƨ1�6��D�0 s��YHߧeͧ�^�bih��.����]��B\d�K�,����|ͻsS�t�le�����<x����V���Ɔ0t�X,:=����=K�Tm{��2��Ɇ!�%�p��/�����Y���5n9��f6b�����:�^�$�w���ߚo
���L�T���
�0���x5C��j��3ë��ʍ�K�6!�����,�Ⅽ�j	�]��!��3����DЄ�a�Pxo�`2�{T~�ش�����qD�d}���g`09(FaD�b�씜ˈt{G.���xǪ�� B�(	����a�8�ک_��6|M8�� !�sg#���=�n�7��Y�q���dϴ3Z%�nص���;��orBh�;��f'G{��R�}]9�6��,�=("�{M( �F�:�5��%nB��ߕ2���;Z����T�:i�n��7t�Re�Я+"�{��L��I�%V������Sg�h���X"Q����FD?�ʤ����3�(��"�?�-��mCja]1)���\�z��s��9��P����C��y��Yw��"��wg�e�^�o<2�����}xd�:�9��)�-(/E���m������D��,3ؤ6��S�)�C���4tx�&[��7�cr���M��M(��ӷ����G�ZR�U)�m�{vp>��4g���'����{�?�/A�I�`�-@}j�J};h��	�E�TT����vJ��zjpҀ �az��&[����Yo�0??Yx"O����x�}Λ�j?A��t��b����Y���@b�nYl�q�]�b!�h@�$���r���w����m.��"[��@&����h�g�/�S���È�@�����a� L������I��ӗ%�=�/v!�-���jpr�v>&T�7��x��j�I�Vx��I����.b��d��aXH�oc&�uu˥���1 .�NrSS�`�Q�xEjM)����A1��:q���HUL<�o+\���+���O����+���Z Wp�I�8���l��j�/�Ȏ�V�0ƛ8�~��SA��>�gH]>�Ǿ��P��u��t�Y��Dd�MW�C�t�4����0�`W���|V�9��8�=�<T#n��K�Al��47.���Y"��C}� �^z��Q����K?ɞ�2":�\b����7t��T����c��E�қ�r�����r�&��j�@���ˣw��t����z��p}���S��Rš��yeP̃����M5ip!9=ļ��V�IѢ������"�&C�nL�V����e���Jy��sl<[S�:��Y�P<K�۵2������w�PRǴ�Q���66ԓ�=D���o#L#�Ƒl��̇��4W�^��d�x�&E�H��z��G-#�6ze��<+��������K+���
�|�c����~X#]Ђ�AiE����A�����B�~� ��%�}�� ^>��`f����/�Лp��.{�F g�E:o�����n�u�e�jo(h"ev�!s���ˎ�� sBm:s?���:��|�d�E��Ϲ������D�1��K/��s��!z~_��E��+�ڔ�$�"��%��"t3H�<z��fZѯ3~�7�����!�:����3�u�M�R6ày�hΜ��:��x��q�˕u|��fD��P�� 2A�/�҄�Ġj���k_����� z�ةNg�Jvk!{}Z=���7j��1�q骖MTŒN^��z�'ǆ�gV�h�0(�?a��MK�L�KB4 C7�7�� ��������?�U(���<8�?���9�޻���s`Ö�=��{��A����	�[t����{����������I�S���ڤ��hgY����^~��䱁�w��{��?���G�peȦ"�vt|7,�
����oGbFB�S�Y��?�$4��g�*[◴UȆ�3�T��`|�D���?r����~���+A�[���6��%T��C�>�"+P���P�:�����Lѵv>?�h�;��3D���7�/�nd�W�
���Rm���٥ [mͰ��L�=YNV62u�x�%�%�!*��T��{Q;0�W(��wu"]2s=��:�g8����O��D`���A&�r
���+ϛ?���w�U@P�{�0Ղ��<MZ��=
YmV�
_|S�7�}�2�@�y�Z�$0�,�j����?BD!f����p���'��[;�ω�EMl~+F�����뎿G
=E��ZL��E�|g2!�KL8�u�u��!����Ks��q�5�]:�:|o��Q��w^�"�W蝳�:	'Ӏ%c!@#l��>Pn�2W��|�;ԒY�M���=I;
b�Fq�κW��{�l|�2�B�B44�~�}diFb�R.��ۨ\����r��d�W�����yFM:.c��$��v�ٚk�P��P�݀k
����c�A���
[^�.i߂=�nB�j ���K�r��H1��V�J�'jF���M�O:��b���j��'wL��ɞ��8��n�O�	�Yݽ.N�&K�ʼ�c�o����櫪v^�lBD���ؤ�2(P��7�ۤ���)��)O( ��,*�W
���_�n"��8D���+g�R��yK�ycg��#�Ѥm���<(���t���7Q�W���ߤy�r!"�SJ�,�Yƌ����(�'��%ڼ�KjRW��{�)�Sܽ�``��g}5"oH��9"o=o�-t�4�Ey�B+E��7�%^8=���d?@AҐ=/�<��G�rH�X��sY��+�r��2Nj��|��y���B�<'���#@I���̧s��ސ���1���P���6�'�,C%!�la�w�d�^�LQ�u�{){($[d�w�A�){v3�΄c���5����������{��<��>���b����ݗr��,�6�o�V�_��x�W� �Wo�B��|� �,���,���E��>{��)�������U�د<���A����g��o@jV��������L��勹��4�����+�bO�5)A7|��{����Z�l���SB)~~fȞ"��uq_"N�Ӿ��Y�z��۩[g]�)e�����\��;�����n��'[G�E����L��q�j�*���+�0�N��i���R�[|�15�bs.#�:sH3D+du���=�[ý�,`�#�kNs�s���!mkk�|�|�����Y�����ݡW�u�yk� yQ�� �K�����g�j���T�龏Ӓ��	���A^�Q<_9�������j0�~�S�=���PpzF���[�(�َ���g�ޱ����9K��	�ui��q��:��1]��*�n�P����5y�D�꫙�:���ө�	%��_h�.QQ�BY~�@4�f'��sG�L*����g?|=��;BgR}����R���9��7��PR�QhRK�9_O��l�ݝ�ʵ����S��M]d�*��K��]5!ho?�P�?]�x�f�B���=�K:�Q�.�]*�ۇiŗD;E��
us���&[��.rt!x�Tw��X~��� ���3�\-����g�ZWf]��*�x��.Y�L��׻���X}K(��d;�x�4��J�J7jϗ)Xߪ�[t ������з��'%��[�_��0�_����a���Օ)A��7����k�Vۋ������?�S�:I�'p�Ǡiς(Z���4W�v��l�Չ�%�5���n�:��kX��W��޵x9;Z�� �N9=�����Y5ߛ_�
�H=�@�8�ṵ��E]�V;�C��+�=(3`2��QU2\�U��ZR�P��1q�J;�c츅D����θc��iXP�W�s���5�nݽof�'yo�q�e��9Z��k�]'����5%6�#�_3����N��>TyL=L/���tp?r�_�U��1t�$��#���O܊QN3���漙\��qO{a�w��|������dv�}hRI���G@���`LJ�=�+��G��t��FP��^c�f�����w�W�/&/�(��o;�4�\��:�Y�4@~C!�.�¶X\Z�x>��*�ez�&]��mkk��N���D��ݹ$�4a�zL��S�}���0"���X�x휗�]p�����j�n�ؽ����+F�ka���ΙΥ�j�k޶�����)le��;O�3�39?5��b^�T�ܝ����:S1�.حH<�y\X�f��N��| �>[��N��5X�\0�Z��c�˟��M,��[I�ʕ| ���?�X�ң9i۵UEԓ��R�_l����FdR���7���q�N�Gk�u(���[��t��̙��
ʪOF%Ǿ@햄��1��zQ�ϠP}�����S>�%�������}�������JJ������������h��W�G�4?�ԋ�bKfY_$6���D΋[�����Ӎ��%P��x7R�3�ߙI�q2��~Rj~Ys@;OM��a>�p`#*�W�ʨ�"�"dxy�oS�3�o���������HbQ�Q���7׺��㶇�^N�j�Nѳ�ŊY-"�
��Ѵ��uLԒ�2r�A�|ڂo64�U��*UϾ�/���C`+�g�)��V�,C(��S������ԇ{�O�HyG[a�z7�K*h8���X\X)]�4]%9i�KK@rY$�n�S"��$�y�������ɇ�r��c|w��w\<J�b����9��D�y\�!�p�>D�/�ߏ[F�zg�Bi��-T�[�Ϗ����0v95ȏז����߉��22��!��Ɵ[w ���$���ei���;�D�+k�Uhk�{���aD���]5Ǌ�T�)Ej�0�|��7}����a�B��G	\ǽo��?{тf=��e��k�B4���/%:�����]/�:����^/{n��n��;d�}�ޘ�zx���m�����s�S�j���D|�!�7:��o�K�\Xe�j��Qi<"�OMEk���O�)r�7h:LQ3�A6.�C�����w=�p�G��&�:�15�n��2����A^��ִ��U�3�vڭ�Bbd#i}u�(�p+ަK�+L���^����؎�ʣPL�H��}��&�p>�s�-��0�#K��&��A�}�r	�\wp����EGBfuuk^5��aOp��F�v��
�j������� �i,YWϝ��&+�	X�L�3;Xf�� P��V� ~W:g�q��"\?9�.�b�Bdi�g�mZM�&���q��,4�J7�C/�v�ߑ�U</m|�`W:@p��Z�=~��A4�q�>��489��������9y ���m����o�EL`s�]�J8���E���v�<��iY~�$�2G�ה�4gŊ�O�"�uӇwÛ���FtKo�t�@ ]�:{V/sI��j!`f�x��	}Yr�tI����GL�J�5�1��b�A�3��2�q�LA�fj�V�����$�y�Va�)b)g�9��s�/��Y�vV�#O����G����p��-/ ���g��=�����!��+p;���_n&B�L��� Px ����^Qd��D3%:o����ʿB)p�]���>����W������Y�=7�����8q�R�(}���/^S�9XT���w���^G��eS[MJ�YhN�Y��/�&�j�GY���L�l�_r.���q��aE*NQ|DݛZT�����kq�bS x��L�x��G4d3�hBX��5�W#�mG{hd�^����݃��U��q��g�ҏ�Z(X/~jN��KwXsZ����1�^������.GE��t(����/b$����t�S^{�!�ğ	q��ή�o����8��)�=Ŵ�K#nJ@�+��#ݫ�Ҷ�p�#�F��Q|f��Ӣ��߸ܴ�r�Q����JSx��k�;6�@+�h����bs2^�^���@�N|����'L���USG���)��%�߆[�E�s�3�UW��+;�x���>lk<�EǛ�_Z�~�ܢ%dSK$4o??��[�lN��&�sW�ab�2[װ@Ap�*��3�<���d`/;׬l��[�{<��~��l��t}W��6Ԏ�8&�->�H�x.��k����~�m��26U�hN��}��`{�x0�O����E�,�xᶃW�%&OA
5���3h��0��=��B��"�o�ϓ{I���Wɘ^��/����7�W��cf ���a� NP�/V
�+��WT��co%������6�����6� �ͤ3����=����ྖB�Uy�
U�3*���VR:~L�;0~�,�� ����Ks2t8p���:f�7yD��N���R��\���P���0��Ei��CJ�n�F�z:�X'&���/nE�P�䏌���[*u�/W�*d�a	.�(1u>��RVMqL6������<?<����A�7���K&����%s�V�cI�;�h���~r楪�1V���R�q�?�EG�o��+��C��X.�\R���.R�1�"�إ���Z�����<��釚_)/l��L)���|���V���˭�h!֜�,��ܫrx��n�"��dw���J�����<������8��Gw�"��c�)ѐ{w��1W��|X��,�U�Ӆ8�lA�� ��<D0v?�o�m��1T?^�� �%�Q�ư�B�H��PIC=�Q}9�n�X�\'g�d:>���:{X��:��7��I.8�c����k��Z���ά�h�D�8��E�j�;i/h� u}w�[$�o���;n�H�V�̕��w�X��J����CܛE��9 ظ�j#0���C���B��b�����ze��Ũ�LXn�:LC�Ǳ��4˘��鹯�羨��(��}�X���,�D"b ������5��)����r�s8��{��OOѿP���<�Ji*�_�?��kq#oů�C�o��O5r�j��Db�XI�7�$H^9�@��C�5?��	Jl��R�\I��J�[���}w�'WN�@�11`+/�w�:�lGm7t ��ەm��/7�+#=[��z�P��t~���h�N�{�1<r�p[6� ��R�[���	yM
�r�E��r��#���|�Dc�vo h';Ҙ���8%osȪx��|ɋ��4�o�Qq~��
��bpp�L�'�$F]�6���c�V �g�P8D_���?�����܌�G�11�y�$W;ܵLC��f����a.��z-�z�u�
���2H�h`N�C 6og���̈́�>�A~-n�T,y�t��ua����4��zu�2'< �G��}��-�Zj�4��ӾN��_�~
�\*����a���_hך�@��{�.T����'jOj-�ݏ�L�Q�qôn���[������4�Mj=x���MoE%5fA�CS�W3���Ve�Z#��E��P*��[�Yo��+�������;e@G��"{�ݗ��\��u�횩����MTj^��+��w����yU3�W���U���W���8לF�í�2�u��!n�o��
fM�"�N�z���ު�F����%��=���4��ۖ���l���O�b���}��I6����̕��]|�WJ��}��46+_FS�����:YLq���)W�����G>���e@�������jh��7�f�%ڻ��s3��^qƃ�0[U�e����ǪL��^��-���n>hH���~��=]���n�C�R1 �'�@��r�_&�vwO<�-ޑ�|��')���75|̱��v���p�'�z���$�b��'�X�x�	���"���sL�?9 :�m~��\K,��V�l�8�
�;��[�N���7�H�ўk���w�����2+#KU��k���Ƒ�*{�<�!׍����P��b����3���d�q���N��d�k1:{a�|�@��6�V1:�$���d�Bc���;�$��C�'v�
��>\b�r�mf�&�㦜<�Os��f�������֭W����t��>_�1���8�j�`��C�Y}O�.��߬�P��/ �^鎼w�����,ؤ���k!a���D� t�� �f�:?X�E9u�Q	���i-�9�"��|^�����V��i�d5��!zY�b[鶽�G���C�CB�0�}͙�g!: a�����H��@"�����lF\(�NM|�,��k�WŻo�g��b�}�Tq��](�lų��'�m�����榑��X�~gK)��Z_���q]��U����7�J���J�+�ଣ��6{(�ڍ�1�<�6}�������@�v̢d47�B�*a5��w�}*џ
���w|v�g�#�J̲��b�A�m}�(��w~R}��B�v��U3��	
��"s�og� ;}��pX�����I�i%	�͏�y�T�J8�#�FF���uhۖ"
��o������8���W��-6^>�/[���k;�Z��F��R����=�j�bï�գ����8����5"�������L�߮MǇ�%&�Ϫ�ȿحa��R�d�����Z  �	�]0���id)xu�����H�k��
�Y�)�-t�6j[=~MS� "�X~�fY���I�`J��#���i)q�+���J���5j3(���SW�o����P�{@3Zgb}�����i��/����E�ŋ��J����Y,�P��f�Ќg�!�$�q���m��\A�8���t�9�a�7A�	�Zf��-0�o��k&|+ii��vpr�O�� �J]� ҹW���mwN렦�u��n��´c���s� kzh	T��(2���;�&I~Y�]�G�_�א:����B]�� k���"H�r���X�x�d|�<� ��a�|�grUn�Oo��/a�@;l�0V�A��k�7_������Ҡsȩ6��D�]�l]5G�j��e��ۏ�&��!�\�9�%�b���������ǥ�F���=Ei���f��H8�gx�z�s�3s}��/�w����d{X�q7�L(�V���}�u�bL�T��R?�Y��U��'G�IJyZ��Y�?6�up�Q����7ҽǡO���h�M�0�%�KVXN����}��{	:B�s��R��T�nvxf����/�L|��؄����׉eT�%�����N������/�Kn����Q��o��:7F��-�MO�.H4�s�]�r�|�Y��>�[�x�2Xĝ�u��
}�g��,�a�� X��+:!����dMB3�����Gn%s�j��t���0�� ����m	{�tM�6߀�UmQ�-}-s^���\m)_��7� �x��-�Z�j� ���F���]�yf���(�8oA�i�9��f.�������3ac{�܈�t����8k�ݯ�u��4��=�~����}�39 ��{��7\��E��	t�9�W��._@��hjM�A�4�D8�m��Ղ7���w�	�߉xu�����Hk�Wդ��]��Z\���%v~e��{>_���~6�`��T�Ԗ<���£��j,]T؞(�`��Ql�8I�z���ʘ��a7�/�wE����B$�'q��^0�G���P�cq-k�|_�ҽ�����몿5~���YC��*S&�%�h�U���7ԊT�V<����t�����x��-�|�Q-�e|�`^���4�]�D=�۹q�٬��;�4�Ӧm�d�EC����<k���� ���VX�Q��w��a�k���	�z��@ܩm��נb��68��Q̲ʃ�#��㭣q��[~��_��%�����G�~ �Ӓ�ZFof#$Ҿ�b��?���1��^���;���=����+���1���Ѱ���9��>8\����`�,�E\���sfu��P��%��z:����,�I�Y-���
�.bS�U�(П��o�Wc�WS<�[i��-���fcX0��ee�&\*�(��r���@�NS���%hCr~L+VJ|�}�v�{&X7Vۆ4yA��Y�L���E1)�]\w� ���M16-i�Y\@m��9�	NsH��7�|�q�����`���1�/�v4�[Â�o�h����AO�4'I�_�$'����}�6�Åu��!�i���>�E@g'l�W�i��S��@Kդt��K���R��W�������ԝ�G6 �٘s���Ř��@�^p��22�.�O6�M��|H���}��<��#@s��˞�ʑ+uY.ʋ��U�k.7���f��}Y��vS��V�s�&�{#w{�S��m�*�c8Ӈb��I�_�nV�|'5WRϽ���X��K#� ��"�_���ZA�^o��w�K	��z�[���G�O|��Ui�P�Pf��K�����˖F����^�v}��~�2�}��k@�Һ��o�ơ�$�1��A�$Gm�g�P��n�U�F�q]]��4����d�'�*��n���Dp>�f�Ow�Z�(�Ǒ��O�Jϥ�'V�::-Iq�����^�.|�~+ڌ%�U��j+QuzF�����Ֆ(X��m���h��+�8K�+�Ͻ������,N�U9w��-"JiY�h<)b�>�0�.,$�VI�&�e�%���Zۻ����".�6�;	�$�f����ӭe���y7n�������U��,L�em��9e���w��V��+���/�<^Ѧ��i�L����g��y�X%(~�S�%r�^᷈��Q[Gq��1C5>�E�{�;Y.X��xÅs9gU��뚊6��?z���'���R��;J8} �]D�Ė@p_h!B�J�^e`�ؗ8C�<-�Bi>�+����T��N2�z>�/�pbJ�������*�\5�S_��,u���Q;=�V�ӽ6i��:MqA�}�Ʌ=\B�5X[�[1`��Q�/匥�Z���P��2�R��S��aUaj���W/�Ǵu�rЬgT�񡳌ίa�?m�f��MoHOҚ�Ws�Y}'��-@���/;*A����Cz��u~���=��uXUxmTk(����y�t~W�6,�/����J�~��M��w���s�}}3;�?��"w�҄w�-t���Ϫ8�%��{8�uN��TD�`�ëW߆�����������\ɚƾl�,��|ʜ� �XK!vZv��-�1&_y�����b���02:U%���"K�t��������h�P���2H��+���nDۄ�۱�ܙ�t,nJ,]�Z�� ���R����5�c+�S�M��`�*��b�3"��=�����{��;��`g�>��1�r��%�u�/���$tO�#/�Z��%��ML�)J�S��B��-ĳjk�0?��uP�w�ۋ�)p�UЁwǳ`�sD������^��^��Aw$ϴ-N��'\��C�O9Ƚ�7�����U����>�uk��&��I-�k6A�B�m4-R���.�+�<�oM7��fMeH��X�X�ũ	O-� 1���XE�Yt�
��ﴒKO)VJY,|�<�П:3��r�0�:�k�*��G-�|7�Z$�"%�wF�r�E�W�"-N�T�~�;/(�?d�\���\�P+�k���� ��=��6��{��3���
�l�C���?�M����.P8��ٓ����9���?	�/�c���Ջo\
�	Z���."����(�ڋ�\�v+�V�lo�N��Y;�/�y
�F4Q�6�o�� i+Y�������ѧ5v�χ��i������������XvL�Eg����h��So��5�_�tR�!$�Y.���b2;�$-<���u�×�\_|-��s�E헊�/��?���+Ր��1��G�q�_�1Y�V.ۋ5�qw����m�q2������f����p�N�=LL�h�v�C'�?�pRqC�ِ��!5@:����.dHʏ��?P��̄Y�b_P^Mf�ѹ;�Kpϒ��^��3α2"��6�ךv�u&��,џ���/;�g��;zk�:F-�L*#�^�һ���5��6�����N��Qc�۷�2̻m|���J�짒��%V>nBe�p��s;�'�~h)^�8�"�+���`�U'�+(�`�X��Y�,���h�M��_��Qu��g�t��b�����i�K��0̕a%=���a���<��apZ�3�Q�p���֨��A}�qk�}�@\NSD��B�+	����׾�@S�k�ȣai�bӓYT����U"/;����\���پ��ˌǆV��"�tf�N�$���D��ƿ��2�R��rx��t�a.)��/@Ϧ�R���,4+ϑ[<�-�X�Y�\e{���gY��+�b�Ҡ��/���vV%*����&������E��}~i�Z�~�Uي)b���Q�sTJ�~�ZZN�W�~	�wp/SG�wx|�*�؞�ūVa���Y�l
���J�WI�Cn��-����.���dש�ݹ#��v�4x���>���Z�������>�/(���ǩ�%����t�X�╣}[�}:)@iܶ�՛��qw���u�c�
�w��k�4D� �F�j�^�@�Sp��|n�b�Η�i�	'�n�.>њFE�Q��� �~�l�1��G��q�wI,�5�Jҁ:�	R��A&^C�]7N>�f���n���*��l��8�+4���K ��=���R��\ ���4l]�7j�FUN>�I8��w�@4XinLj�v9��K
��u�E
���/��)���ؐ6����?�?`*>(R��e~)d��4J����1�֞Z��y�{��q{d���s�
D@�cBVvq���+`g(>)�OƋ�a���/d����FT��R����ORUٺ[��aߊi���˫��%�d��nEΩmNG�n�>9���k��[)Cq�B�ñ����A��n��[�d9�Aĥ�}~5��V��+<蚽4�φ��̠ȇ�"tutC�=�Q�=�5A^��f����)��F�m�v�R#C�����~�Z�'�����C�~��>��8o�b�b���x�p�n2�W�F���"J��X��z�7ǐf
i��[R�h5k� Q�b��^�Z8���vjH���~�כ\I��.Q��wC��=����^�	uٝTv�'9~U�Uнd~�!,x�x���%FG�p��������'n�aħPh�=�@퀟H����u}tb{��;)��b������Ƨ�?`�#:��eI*v�U��8b���$ݰ�Ϸݟ^�^���4q�ƭ�#��7��"NC����x�-�KU׈��7��O9�	Ol�+���;�[�O��������"	��ۥ)_��L"yy9{-�wj&����"d �Qr��gM���gSx��U���fZ��f}�8�e��Ϭɏ������,H��ѿ�Qy)�!FDZwDiP�w��}$�����KS����)V�CF5������4�����@VmnM0"Ѹ��f(Z���8����0㺑�)�����	r�?j	%+_>�P�	�T��4𴰹�Y8��y�Z�(�����W1?���v���vr�=+�FU��Քͥi0=r�mr厬���X�-�rq�t6p���d٘��g���/w���h��_qB�}*��/2V��;^T�A+���C�
?z��(In����HϬ�!�F��5���? d�|=�/=0)��Qm �L.^�-a��6�Z?wy�e�Ο�_�$]e�mX��a"C��[���������{� �sS	��īA4Ȳ�+�4#/��M�b�������ɣR�Ok���ʳ���STP��_E��Б���8WZg����)!dg�|��(Wȝ����S�l��T��F)�㬾¸#=Âtv��żfD[G����<��j5�^H�OIm�w�*����](�dsB�`A�{�q�W,E*�'���9M��J��ƾW����1�?SgtM(=>���� k
/$��W�����b�c[w��{�퓈�}�c~sLx�)��?�ʯ�la��9��Bsyg޷�sB��5�J���O�;z�c���F�H1����+�ͫ�&$+����5V��>co9�n[:�ݻ�ư��?!�w���y���?��?S��8��ɶ�b.��ZR��UUF�
���ʪ{�2xŅ��I[:ht�=��c�|�g>R
y|%]���.�U��Z�O�-�7?%���tt��sJZ^d��0�pn���_�����泋y�%'�2)N�q�����/Zx?��j�pc�+�������5ӳ�ӫ��
����Ƀ斅Jb�U��Z��ǡٰ;g�N[�֣N{���\)X�ޭ�&��e����4D��T����'�ai��M�8���$ ��p�F���SW�ܼUa����s_�?i�RPqD
!����N�FTzIh��jZ��J5������VD�/ُS�T���jlYz�H<��]>����§�ǁ~���=�R�tׂ��R�������5 )�C�[��ƹI��0���''1���̪85Qk �s�P	 v��� `�9TI'<��t�.g�g0_�Lٽ>'��ktW1�7%Z�*pg7���$�R.���i�פ��D��&C2V|����{dXd�:�YK� �r�G�L��b�$�S⻃(���Y�UDSm\��Y�t��Ts˛�n��@���,_���2L��\��v_�\(��Z$5��J�%�;���d�{@3���2�{~"8���n���x�ůlN1Ν�Nan7�ԿZ�Dۿ���ia7�z�Z�sk>t$G� ��;Ň�JM��2u��0�y�[�����rg)�I�G0q߲�q���"�pCW'�^hLl����-U3���в�u���`!�q��#�Р�1�q%u�\a/̬+�`���}g�W��~��vM�
Ӝo~�bH'������}��'}�tZ�ZJ���G�����������߹ �\��ǌ��J�zy��pj��dU�;t6�e�XR��aP��(C��^v}�#z�J�B4�]$U��ER��U��\  /�x!8oI��$�8o�e�ߍ.He|Kǌۓm�8!�܊��9���kl�@+o���ZsU�U�9����:�<7�Y+����s��v���w�����0�\����SN��8�S#�ߦ��~�n�v�F�w����0y�f��%F�����ž�d?N
RA���NF2�q��(6S�l:Kf���;P3���B�E������Jj�8$��A�m��:�-F�U�yw̸/�.��$W�C(�-I�L�\�:I �*X7Ø:���GJ�������;<�9�2�`c=wD݂����#�(	N�\�;�즺�?ϸ�'�ߋ���l\%�(F�[��m۟���I�<E����M�YXP�RK[���)���h�[T%���E��S�D�4����G��MҾ����yn��Җ�)-������a�8�<��w��0MzA��i��N�R]D�1�����?(�^J��p��\�"�7J%�N������	Ks�c��
�j ��[p^�_:����m����c-�D���N�oXx�Dm�i�0{���S�;ǂ����~^�'�B�Y����k�PO�;I?���ƪ���rŮ�C����q*0}�(��K�&B�)ah�dݼnBu����BY��(�bH�f���E.am�nƘ�ֽ�e֪���Y+Ivh�^ ���7���T�9�cD���o�F��tp˳l�����L'��z���4�'��#0�����̵�d�-;_֥j`�l]���J#�i�t�n;C�E��[�~T���X��$n�J]i�z'�|��$a��<ױB�t{p78�����������hT�G0�GUO�n::?t�Z�e��9Z���skP���]��X���Q� U��F_v�g�̕}0���pMFw�|�7��dc�k��b�pO5����놣�Zw�8_�$��a7=�lf��_��ӌ��hʛ괶����&�ٍ�)kB��)��3��P�M*C�f ]7����no l �� Qp���kt����/�+xЛa�a��5+�}6�7G���j������vG��݂��ujF�wRs���E�}�$�&HѶ���:�����+�o�F�I��.��C���Ͳ�m�R��M/��!�_�%P���8/;��� L���t ��F����0��/L�s��.[��b7��5--L���9�U�gQ9�u��G�v&�%�v��l�av�@��ܲ�tJ�t5x|R�h;B3���H�(�x���q=2n�L��[џ���ͫb�<�(}R򐻐28�����[|5��?�&<z�$F��uGh32�����U�d@"`�H�T�����W�F{WRM����ӯG��*30�Nv.��/Z����B	�'v��'�5K_,��|��O�wcӟ�y��r�g��%������t�ٳ���E����F�F`������G` �Ϥ���Mf��x�ڬ��QE��U��S��e�$�/�g׊/�^�!�L��<���9+����M�ܔ�v����݈Ɓ��ע�?�8��0�S��������}4���}�q��Gx��rZN���#�h5�h��!��N�^�mW��|�����B<pp�)�\�`��������I���
E��,��,Ue�l� ��ౌ�H�5�7]klS
�C�.��N�����2o��Tc�~A�2����d�dE�CÏ�Z=Qԇ��M\��	5N��p�����E��xr���׳����m��<�AM���_@E�/t%�G73���
�+��y����j��o�����LMѣ���T#�F_B�����p��4~��%���$�8�T�D�{e�%�zS�<,�{k�f�7,��j����^xa:P�i�0 4�3$x��;�9�~�]b���5�~��s�S�/�!�}M��%7�ɨWo�� ��UzK�t�n��Q�F�L�_�iNo����z�P����e;��7e�B��3[Yp�X[��/��R͊���v���\�rC"21�Zr�n�<Kd���������#cT�"�7��@���t�xϭ~�A��[��i������ǁ^M
ZF��Y��$�f�/�A��cj��$���/_���+3�����|�3|�����mʏ$6�<���	:h&=�xT!xG?34���� �{?��:�ngc�.��VCW7*����y~���TH0t�D=����̊�����Z��X�>�g�У���"UF{w��?9�8)����VY8�{��kO(Ⱦ{�n�R
��]��������?��bWu����8����� ����~��lxGo�͟��HgP$/�5#X���L6n�gO�Wh�R���2&�Ѷ`�&wV��#xI懼{����t��ݘ.�8��𘙮{�~=)�z��-�$���e�^B�-h�xqU�W�"�2��`jn=�e5*~��T%���p����g�ڢ>��!�-�:DmR�.�Ա}˙ɵ��#l��|�1�/.����ɀ�j�q�״re����"өDt���Cbk���>Ѭ�V����TNe�
��������@V��ѧk|(*/���D��
-irYF����>�s[,�V�C��7+g�*�o���m�W>�?�M'����P��G�Ru�N�G3%�Z�j�k�Ó����U?L�p�pl����0Ӌ}|����,��ro�����P?*�'�^������T�g�I�.앙�eP(�=4�e��B2�[�ݮŖ�`>kL].�o���3����=bp���r6�-vDr�5y�������11\o�g���:�������gEփ]���G�(�Q��5*';^�6L���+��ǧzJ��doc����P�&��j^��A�`ݟ7LL���̗�Z�#=��co��2yi{����$�	�p2|7��=�O��M���+e@��>�=o��3nd$���SO����n-E�穖��|z.+mwK�0;k�כ��A��q[�S��G�QMY�5"� ��oL*l���}�� ���U���L=� T�.��T��%�FM��b!{�N�G/�o�tf�6�`wLO��m�#&̬?�_l�����}O�*XͲ�ۑ/>%�����A�iS����+�^��}�����M����Ax�Φ̡֗�+��0Og,�@6�Lק�Yb��>Ϳc�?��:�dW�L�~��RA��n��i�����Ϋ|
�Y��!i�I���Z~@�����	*2���x�����Qo�f��M�i�h����f�*A����CkZ�����I�!D�,�v�u�ϯQl�k�������ݦ\f��Ӭ��.xRd�k��n��Q�{��oEQ0Z�Ұ�Y���w;�3鳩�t�%m���98 ������ �� ���R~�i S�3bBA��Ag�3�0k)�b�D;{� g��/z��"6�c�����t�f�ͬj\���N���Qc�Z�������e��-t�aj48�\5$��s�m�×�H�[�ǤR����)r�g���_^G������13H�}X��=A�?\�~�9:xp̰�e�Km_�Rz��Z4O�~@�:��7�P.j�/BI���&
����3R���`��LS�����'��Zg���9J�u���2�ד��vPۆS�a��h�1*:�������З���g��S�ߞk?R����z��|,��O�3�Y����x�j@d��t�Ϣ�;�v�i={n�H�VVZe�9�C$4��7�����F15�w��=w#3�<4l{��s?S��nUh��N9=������6�[|��R/��׊fY�U��؅r��bc �B[�H�8��v�9͇��,fJ{�^�K+��WQ��˜�d�]��.AG�śfm��V�{��䪚 n��iErI���6t/��؊ڌ�s�/
*,b��@���Z��g�Z��9� �aJ�4f��h0/����'������#p�i���;r�j��A���-�T�Y.`�,�J�i^��8n	p��&�Lo,tq�I�"��D9�)���o����k�/J��H� ��!av2L��>�>��a�m���na�!c[��ԍ[�����⧱�q�-��n4t���}����X���e_�,a�6 J'ˉj�Q��L1���u.���?��lY���r-:4�߷A�����W�	u���IC�4y�e���	�\Ĺ���v���/�U
�Z~���-���S^`E\U���z����B֮ь��gddd`�T�;�DG�F���BU�{��DrD��c�I�U���\�%�>�1�/�E�������n��#�QuH�=�����;��nfA�;o&|���9�wY�Q�qqJ���8m{�;zL��@Xv��5��_\3��Z�d��&¿z��a����s%����#ӿ뢡U���i{���2�I@_��m�+݂';t��w`�_L- �z�d�w�P{�Q��r_��d�/�:�E��yR+y�",eC�f�|� B��z;��t,n6|��]S���4�|{Jнm~_i���ݍ��������H$��iO����u9:�!۴�A�N��w�W���ۨ�P��}�o�}�h���
_�X���q�]�n�
kjEsHT��V�����s����o�O�%������x�WG�}�r5d�n
3����ǥ��1�����@q��wǁ��p�˲N�!I6�}w���;�i���������ֽ�L���>�ӊS
[x�my�i��kpd��T����b�h��A���5�v�W�N��Y�2V2 ѐX\{�l�����s# � Lͻ7*��K����4�ݻ���,����/qgk�����AU)JI�=�Vq�<w�-��YZZ�j����X_U3U������T%bLT��� 	b�{��߽������t?O���w�������Z��ۉ����F�_!����F��ڋ D�5�<�K큄y������A�k�X�:� ��}�o��L�X� 	^��=���ܝ~���v��y�����?�m��a!.�s���D��(
s����!�����B��ﳣ���^m���ҁ���.�cT��Xt�W�d�uo1h��{'	�b�=Z��ք.�zz�p�����=^��6e�dɗ����x����n��:�R;xe�7,���\�^Z<���R��iٕ�%���:ۄܐE=\W'4��A؜�9kO8���ia�:�p��+���X�)�-Ġ�>V;5���:�2�Ǟ��������g�5�����(oa[�2�e������iUdOXpZ����c��?Χ��F���������,�??+:ڀ�$}� (��Pva��2����d� ����=�1w>ӱ^��Q��T_k��qfư��Q�@�h(S����󹎽�p_��bnB��d��qk��#�]��s�^*;F9��`�e���]�b����Rƚ�̌�r�����{�Sb�X��ر�4�)d����7v3W�n4����W��C-wiIII}�+�7�\8��m����>�OG��0x3�������������6����e�|u�T�q���H�9�̓��<���~�lHV#��n��(!��p��{	E���D�L߸ޒR�,2zYY�"�������-��b[�4��)�,�$x_��  |����S�+���+�M��c2��g��d:^��lG:��Sښͥ���q�tSPЦ�YGB��z�O��ɣ���w�F:w��;\ͅ7rWF���_ygX�AB���9l��h�[��6ԣ����\����2�f���y��~�!GW��;>*e�F�=��P͌O,��y��O���
�����2��|�^ ll���q��+�������,�p� KN/1����O-�s}�.�>�幫��긄y�d{Me���A�@�#�1I%���AGW3e$w�82&�,�k��~T��?J"v(���;�����>�����5,�?;*_w�WE{�����US����d9U`�F��7��P�� �sj�G���S��X|�>.ף�����o"�9{����J�8	"@'Uh�j�d�Hu���
&b��k�Y,2?b:�vu���qM8�
�4bG�>[���v)�[/��Z�C��=N}-�ɔ��˭��n��˼�_#��!��&� >ɭ?[o;��|6�`pں��v�ؔ\����<z��(�thx�YH��06�&�hg˩���E��2a�?t~&�*o,��Si}�n��o�F��~�����%-����Y講5Np�qH 6샗��G��X�[�ŕ���|�R���塯��		O	�e�|]}��`g�Y�"�^=�l׌λ*Y)96c20���8g�L&����x�.����3ؾ0���n��k �p�:���t�i��y0W�=�=�z`�'�[^�sSxxԃ�4�����I��KR��O�D��C��^X�����(;v����G7�*���;s6[j���%�zi�b$�l뭴�����lӥ1�4���˱�\O����7�/�jv��ߗn~�N�H�x���Ɂ/���P�󏣱�j(��ҙڢ*�K{������4o<��hkˡR\����|r��M�.'����P�.��/�/6P���dJ=��lJ?�~�~����''vI����E���m���ɩ3�=������]1�r�p��;�U?���p�lH&����ʓ�7n}�w$��'FrAK��L��2�/M"y���)���[����-���w����ݨPi8zSck}{*�d��c0�iq����>i����o��&���Cg&n��|8�W ��rՎ]eiBXq�8��q\˟���"֗���)y�]z����S��*��]�a�!�Z �� N������;�#w�_|c�a�(^A���E�'��,���]�?��ϋ,J���� +���h�#ꨨ��8�| ��;sՊ�ɝ�t���jAה����P->8#V��Sڵ�8�X.v�g^��*�[��T����j�V���S�Z���[Xq~=�Zx�ұƖ��7c# )Kuԉ����M�]��;�U� qҺrXm��O��l���w�|��1��cx�GBZ[|8��Ҳ��������'º���0N���E_.���k�s��� ���Q�{��*�"�t)�X�>�8z���Uaڭ+w��3-<�s"����J�v9g�ɜ"[�F���y+|Nq���d�����"��Â������z�
��WB�� R����Y���^�#��{r����Z��X�����	w����T��?�s"�����^B�BZO�8k�� ���^�c�-�
�=��~N�t��@���˲����S��#X�eo�8��9��O�i{�v���������i��:B��
�e�#����6UW5� h1��_��G����?w�}�|�u���\������{�Oqw��A"���R�p9�/�C��A��2B�|?��z!z���H��O��%l��qe��	ݚw���	w��9�r�i���'j�q�5�|ŨKK��!��	��e}��G#Wv��syj�u�����W'�݁�'?�Y��d>fIa�ё>��X	v�8�fL�oon��
WsW�9g��h'h�Nhzt|�&CN|c`�p�)�l�0t�
ߞb�0]t]��M7����z!w!��d!v�ۺs���j���
<�r{)-�vx���vx���h3�^6���Jis�뷉. �`Ｖd���VZ1���31��^�_���M�;V�4��L#IWӦ���Q�C��}�2��"�؏`�is���_�S��[��by�7��-ܛ�	c�;�G�ƌ�:%Q��L�^^sC,����s�, �V����:���oy12~��A�7�B7V#��J�l��5n�o�.����r�狱5��:��Ư������jG*��8�uٹ�%y<X���Y9ኸ8Ԑ:]�}�ϛ�^�ѽ@Io8�S�4��A.ղ�؜��&�Į�vpK�F�s�7�F�nXTx�?q�%�װ;OOr�{S��ⲉ��ð<>�*�9
\����B��	J[L���m���L�&��*"f�sV'�T���6�/�
_}Db�}��VUN�yNZ_�%�+�R�x��֬b���-h�b������`%�^�c�ܫhO�׵���)���d��j=<�v�����K�h=��7����TV���E�+))9,�:R���y{��������~������2l�>��Z�9�Y~k������t ;���!��#�%�h5p4D�T���8�gl�ٙ����N�8!��s�c(l�"�,휺�kw�鋋�������3�Y������f��\�@�fu_{��g�A��C�1Ym���������B���c��|�����&���F���+��;�&f�\��?<^e�i�ⓚ��۬-�`&E�Z{�o�~T ���L�S������S����'?g�_�Z�S�ۦ���!�����e�y��}n�E���BKwX��\����P�A��Om�>�[�;���[u���$I�����ŋ��,�	.����lLE�v���쵍�����	��\ :�\sssۘi�S�y�pIke�D!�<����[�񹹹��G=S�Tg��X�
^�A��u����I#��,�`�j���(���d�Oie���lz�=�j��9vi���K�%�~o�⟃�&_ow�+ª�d�$�p�4�\�$e]\���g���R2Z����tw�@l�on�E��+i�/��iF��� ƭ������X�Z��\�-��1⑞~��-�Zkķh����~j�F��'S�-B�H�+g����3����%�w4���7���	+ȧ��S}\-�1D���Ç�i�+��2��SF얞���vY�g���ۚ��^֕Dj^B��P�!����r�_��B"��?H�U|�Iݸ1�b��Tܜ4ӓ��/���0#=�h�q�;͓�	�?6b���o�:U�������X��� �ֆ�
��/b<h��3ҍ?�\��;eͰ�(�����jr��̱2��{35f��Փ���p���r�������D]��-�Ӽ*�(g�ջU#)7���0|x{�h��6Q����u��ߘcm�[W:����F�����`lVIcݡӏ^�ӳ��_�wz=�ɰ*�*&$�����{H�A׼\K�h]����!�>����:�!��`�uQ����X�G�{u=�'�݄�:}\^'yM
'6zM�G�������S�q�d*��%]l��{](�%n��Y{"%19����/ɨe�Ú����e�Y�-�]Z�'wS�Ug[����Ud��Z�("���t�i���Bs�aU�{ǫ;���Cpȹ��8���)&U?��%Zٻ`'���voXU^C��Y�{m��k*���ۜt:��~�#=�E-��[�#ݎ�E��9l�a{W(�6��m�Q`B�n�CzUA��?փ��kuV%�v�!�W�V���u�{r.e�y�-��Ku���#�x��T�涗i���1Xo@�Ź��;�Εu�5Ӥ��?$U��3������켎�X�Q��g5��UN��d�/�J�I��e3��w1---ٴ!��0�L�*�R�`�~bZ�Ͼ}��D 6� `���������?O���h�ߥ	_	�OtJ���2��g�k�K9~��ϟ>���BשKP�N�� CS=/��}�.k�>?�u�&�ㄺ���]^s��-{�^�$7D�|�o�����${�������1o]5���$����,N���V��Lkxñ3��㠙&�>�#�]F[m�.su��X%�2Aǖ!6ױڈ����k�>./��v�&����'��yudx����3/Յ�ad��;������5uكx�`�| X
��+J����C���~�BJOs.�_�ܭ$�H.[Lȋ�l�?��q���1���<g3�^~�?2T���i�>��ųg_��O�|��z��!��.`� �j�+;\�7O�V����6���@��Ψ��d��+ŷ�O�����2����M��13<��)��aR�CEƀ��t*�<_��m�W�zW|�v�D���BvN\<������z~^eY�z�ZW
1L��u�Vj��@����������V��Mci]�AAR�H������:==]0�+������mb�M+ۢQ�8��a�(�O��6@ݣ1���:,�8��)��-�����t1k�7ܥ�WK�����n�65�}�E:������h�ϫv^�����{d�F���,����ÏW�����H˜�;����c��U]�	���O�e Q7@�� QDR�<�S�MV��,k�wB��d=�����Y�=�E%����FSKS�k_-/�%��6�ɤ5��S�H�MuN|����|�����!0��{��ZU�u2���I�!�3b2Y<žy�}	�����cAnkC��&��cH���ߖ�W�9��.�?m\�ڳu���r9P�i�fk�Z�-����~1��d1��j{����]���p���p���6:��S^�D+��ݒ�б����{��O��h&],�=`��e�������QK�$�����0��-�/^���G-s�q"(���n�e�*v9��[%�`ɕ% <�&q�9�-|����d�e�!�R`oo�� ��Fz�} �C���9�ړ���,��M�&��K̿}<��1��@(�s5g ڨͼ.��Y�ң1���.�d[��A�D'���U����b��N�b�2j��V�S�:n��fs !��J�ΎA�ؔ�"f�Ɖ�^� �j*1� x�P'�L����dwN\^ĪjQq�Dz�2�?����b���QĢ��C�U8�̟n`�E�GU�$_)`��1�>@�>z�|�dJ�8����ß�orϩW�v�/_��\	�����ڗ��a,��p�8"p�8� �y��ɷ7�^�>F���h�%���������yaRQPp���([?茲c�#Z�Ҕ���5�U���H���-�ø���iZ�Q�ZLa�"�*�����^�[��?lGz^���2��fͶRK�����A��ړ����/o��6�!�y�2d�q? �Y�*!H1b��ʡ���Q��6Xn̈����f/��������٘>��d���bhDL�\�+V(~�c�A����l�)�Ox1��҇�}�Պ)2C����L�C_��B;���d��
����w�5��!�yK�+gs�L9ٲ:�j^��%��<qd���o�e�ڠ�O�k�W隞�����4����lW�3{Z�W8��0sb	�(aaa!��MJ:矧ҵm�z�Ё��X�~�V��_�5���*,j�v�a�I�l=�dw^\��%|j1�(;ᩐHk	f��H�򎸌 ���� ���OGF �z�SL�V�s2�F��%�^�'�)wdr��؉�hc��թ̩Z�RѼ�:�� 4�S���>����́zZNWSS3��g�(L�d�=	��ʟdbN� cW�2��w�"��[�ҶZ�D>X��ʁ�aH�[N��9���
M�P�AFp�I��L�#����'�������%�F|]�c]d�u�D8�ɋ}�������Bƞ�K(�.�2����4,�v2��׹��#�t�;:�U��\;��50ssbT���\��5��-�ˎ���M���6�,�-�r�)�/9��C����L��f��<mQ-cZ4�9�]UU0uݡ!@��2:Pl������B��#�9��Kہ���Q�LajGwǷ��aS���ӫ��sW=y�� %h������u&�ɺa�ư�;7�j�cH�p®%[�;��7C�z�C��j�CÑ�!�hރ���%A�.��+ @BY4Ͽ��$�%�s4m!G�ű&ش6c S�pQf��^�tI4�H��UK'!��݁U�*NZG|R�~0�Ҡck����5��ʜ�9y�%[���xN}�xUy��z��R,(Mɲ H Yؐ��t�7�f����~c 羅�Tq���2>��aRUp��[6t��h�J�r���q�e��� @LD�DP�����,�p!���ڠ���J�9��)?��/?�]�g��z��rc�H�W`8���s?�T����;���	��}P���4�x�ܸ��
�_�w0�-��Ѱ��-����:4R�����,�ф,2��A��;8bb<����<T��OcBU��[��E�sǀbbR�*�Ei�
Tb,;yxh�J�	\u�i�l��=�����{qE*��21�4�l����R��
�p�̡�SN���W�er�f�Nej.����[�Q�� =e'm(�(��/�8fP�M�^rSU��~'_��Wo�� o�B[2�V�F�Ou�n��j�^�{[W���s���HREEE�G�e/s�ֹډU�g,����#�!���]�+���yAf��^LƬ2�����d}'È쀏4`�{)݇�1vS�		re[���+K��)�8�lr�G��gwi�|�1�D���M#&�SeW�b�������ܜ6z��ǳ<�z*���Y��(w��h%0����zF��3�^�CZ�}����<�:���Q��˦�K���FxW�AwRG^�R�����.{�c��� l�%�[�C��hӣ��cPǠ@��2�͹�Y��I�;J�"���V7���[\-�0�]�Q�2ѩ)ȉ�a������^�(��jUoT]�M��z���p��j)�1��~�1t�p��U��ͱ�6~��<ǳێ�UKT�O+%�8��^�1V�;���9��%�u�g��R����z4+�cr���(gU qx���)����〉~�|�i���Dm�rv���m�%"�h����yz�#:>#X�D���2X^=���@#l�f_7	�a���ڢ��$[������:��l��?M���~�����k2���6�x��{�s��a��|N������-E���2G&����Xk��Al��b<���Q��*pB�ޙ�6��5`d�uku��DjT]Jt���pě��h]�,������Q]�<�VNi���v$<{#.,��v��sV��/��C��S\>��{ܮ'4�|�xb3}��c�>��o0W��m�d�뤲��l\����uS��Gt��uei�u7�@"�@;-ݼ�Z�� P��ZWmF�}G�0��-_R������ɓe�ā>��W�3��Q~]��؊q}��pf��pEJɀݖ�N8e��Y�)w��2P���Sd�� �B~X�k�ܧ����V�h(.�gƥ��#P.^>�|��Sc	B�*�K~0''ǔ��Km<4ӓ̓��lo�Bi|a�����|3��CJ�k��D�(�����L�qF	{aBZ&��\nKC��m��]k�r����P�kj~N���Ox��%F�op�ޓG4]]]OW&� ��j��3v��Ī�� o�2�t'��t��T@�`=?�l䔘���H@���|�YW��Y�[q;�X��R�w���I�|�J�&y�᧐�#��$z�f���
�Zvء�>\<t����0L�iߚ���21��Ғ*������6�ACgg9�R�L��p���
�V���J��ὐ���#���'B��I�4x	Th�ql: �v�hC��:�OkO>�X\̟���*�M�00�>昬|W�M�^
�`��I
�OK����}w(�]�z�������a��ё�����:���<u~��Cs�R�#NB�nB��lbF�K[��� �|���ccc�����i3��uuex�T��me���*-��ɣ���_=bp��0&Ӏ��bat7�n�6�4�z��+��,0��c9J	!Em�����x�z�7�%��L_վ"����/��䗛�~\E늖1����lud�o~�N%Q�HT/�Y�e���=*y[C]]�z���$�f ؟ZC��m�-��3DI���>�k�\�˵�?�Ȱ�Q�LV��M� �P����3-���n�����{~�+�;�l�>�OR*�A3�;5K�	ҏ�3�NX㽰*-��ޗ��u�ss@�ad�hK �ttGMLxpodi�}r�boAo_�%9�� ���ݎ��������%<���ee�&)0t��e�H���'��=��e�Դ40X��>�(Gh��m1hW�C��e�{C'w�wK�,��z,����su1�v��f�`Tf� ö��-w�NeJZV�ҩҒ�2A�uŅ� �m2�av��`���v�]��ݮGh�f���1�J�8�4���6�ks<z�C��ʀIw�#�R���_�u��3-������`H3*�� �s"��kġ�[����P��!���:�aX;�����l�ܘ�4�
�NR>�����61�ꕢh1I��{-bc�w! ��\�><���ĕ� ��9�SWٱQ�@�>~�:O�v�B�q�]�}�f�X�yN�y?�ȤSh��0�b��)v�0�v�й/ý���]���\�K}�n�w�hF��z��y�+����ҸL{��]_�&��>�l�
헍�)��{Er"2�_؀k��G���QLSn-�Nrv��X�>	�ܖ(�X�8X�'eVL�v�:��Ԭ�cd�qy���b�O*\�I��w��՟Z ¨��X��_E��nd&U���H�S�#�lύKG�I��Re�|[�
L>��
��RCǁБ��X�4���|Q�|h�8%A[(e�=9=;=&KˏH갞X�vc�:vd���T�\�����P�B`3/���D���-LUh�|0Q�z�cu�1E�cX=�z����um�<_�c�HM�&Za]��-���n6���r]T���(@��C�lNN��r� z�.x;O�wԆ��� ݗԧ
����8I�ˊ1��qj�8$"g��-\11QfQĄDd�e����AK���{ºv-�r��=�(�Ġ�'�cjr��
}s�b�e$�v̺��[�S�S5��b�/Fv�v��ckchY
a�;�t�OMH�7϶<�x�n���У�I��x#H$�n�8�j�{S��׮�G����0��Ε��d�zQ<_�֓��p�ߛ�^G����6s'��m������A����������l4��n��;��ݤ^��+�M]��=Ol���lv�ݬ)B(Ö�Z	�H+NPH�X1�;�ףU��
Zg�o�����ٸʈ�X���k�&P�LS��:����hg�K&K�2�R������������]�4��I�m���4{�v��p����;je�+��H���S���_�|�Z�3*��sqqIV	2y��L�r��Ў�! |%�/�����Ȩ���M��,�t %�<�a��h٧O��JL�@��|���r&��,6�%��$�y���l�[�cϠ�o�p��t��'w<O.��d�$�d`=�WO���H~�41�{39�6� �^��I�y[]����'N0z��K�o�����; �
`yh�_V�x��Itj�#)�oi�����V��`G�xX��j���}�HF*yh[��zk���F��+��'In	�D-d
ɘ�2p�ō�]�Ӓ*'�o���k��|��;+��g���Olk�Fͯ����k[�G��?>���! 8��e}?oe� �M--�G��:4����_XW*L��f��S<�@�v�v���A_8��W��P�	��e��� ��nx��R�LM�Gt0��&vJ]��$akK4��V�k	�1�>M>W?�oa,N���ȗ[�$�2��u����t���M`�4�� �s �����k@���Z���D<����	/�1���{�!�z�������<�}���:�
�k��Lqc�g�j*�d��6��v���,��V�-�][�C#��7�h<��c���c_N��qpӽ���� �(.�d�(M/PlG77WJZ.\�ǂBoyc�?!�& � ������ �/�x�̑:��^UOO��w,����/���]������cܛ8f��lr��k�?�P�Kϟ3]��;E�u��S��H#aWkɧ�)�C��ex��_�o�9'�D�E��.�mB_������W���P��ë����ǚ�`H�9м������|}�(�ï���'��Q��H�@�n�2G\��U@��R��7�G=>,�2;kL?@��*�@���D�����y��o��X\��s�sV��/�,&�k�MZ=z�I�=ڌ6Z�K&��FEE��,'�L�??��n0�=�!7X�!�Sq�?�%V��C�	�2�e�{SFv|[��֖DSAoz�S���~[� ��Z\O�y�tf٠Z"�j�c��}��'����������*[�� � �kz���	yVp��� ��M6̈́���s=r�7>)�J �E��������rI���4{��a�!J���ʒ#&������v��\�i�1${~.%=7�XjGl�M��j���C2B�Ɨ7��	��pۂ\]��;lK${Z��k00�ͪ�<~�+>���`��>ȱ/�ol<��N*N2	j��s* lT���j��U�\��Tm�i�~!�$��Aܿ--nvP�4���&z�
!X|��>s6�\[A[�DV���p|xU���L�#1�F���C(<gX��-���{[��W=���(O+K;w7//+I��޴�1��*[wOԄs����~!p�jV^p���PT�x�>* 9877����٧ �X��!�)c`�uvw�2��hĄ����*����^�}�9���T������;���ʠ�?��Q�/Ⱥ�kuh��L`KR�T&��
s}�F<g ����kY ������o��F��SΡ#�R�Z%���j` +¢&:��&� �s��H	X����5ݰF�3��M�Z% ���V���F\ u9�rqʓdW�IZ��%~5��9-x{���-gh��%��?HH�O�\�]<*gv-���|���ͪ�X/x~��^�B<�Ͻ�����<���mll���� �r�ؓ_R���E����".[8�\p�~q �q��U��� p_����������쳏Q^d����/@�U��Ǧ�� ��	wm� tc��fb�K��aaΡ����!1w�ƾNs���A�P	���[�}�	�I�ʲ��__��9�0���@`�'^�~߸���t��^�	�����Հ ��dlߓ��2�M�\j%B/�����[qv�;��*6��A�{��=��i= �%-���:.mr2���+:�s�� ��3������Z��u;7�o�!ۀ�B7&gQ|q�XS��o�7�M����S)�,�=?%iW������3�D,w�1#*��#�s^F����>�5�=������w�H�.��Y�G���gҷ�5��
��5���sf���h<��k}����!K\���|��=�T���t��M$�R�<�4]��+ۜ���P>���k�H�'�(nhh蔄�[�B����t���@�������+U����Wk P����0�Z���������mit��֙++.�Wp�x�P�6`�����6�H��&%�MըY9�	p��.֜�پ�<TL�"{�
X7�!% ے�lv����*�z.���.��w�������E��@�`/��-�u�B*d�3�0XF�Z�A�^|��"T�HRj/$m���7���qJ��G��V����{*��Գ�U��Ҳ¤.`���tH�n� ؓ=�{�Fh	@�$ �B}%!!�ri���.r}@r�.���� �܋�%�����vs���5��>C��7����@:�B��!�	�`o��'�Ç��wq=U�=$m_���@ �N]\����j�?gO��lMc�[_691'uTT�sH����E��F���.���[�VUpp�c�'�<���0d
� ��D�(Jg2����6�&?M�������g�)�`KG�5A��A��ٳg/����۷��� X��1 u�H��}����d��m;���'�A/}��R����g��
(F�#Ե�kK�񡢖}�@C�JGE���@A�~
�3���H``��i��#���< ������҃O���$-V	�rZ�Hls�F����]�+*�K�B��o<�r���'��#��8����9ԅ�����yŵ��r���2k��Z�W%�n�:y����vI	�ӗ3�����}��\�	�(a��ONA ���;!��v��[x z��l�ƎXɞ������������z���Q|��<0i��<�� q�=�tZ��n��ٔY�&�t�sQ��2(�q��SO81陙��*�ku��� ��&/WU%���)8�xZ��y�TAA���}�7�Elz�wh����ń[@ �2@� y�08�z{�˄�o��j!	��{�5�@������i(�B$ʇ��#*
H��υU��> (�xa��h��700���I�u���7p=2o�Qy���EN]��8z�� |�iY��P:r��q���Q_���ߌ�pV@����[�[ǋZ�_g��✿��gq�
�]]u ��^8��vf_ޘ�4{%6ށe�p�s�h SYL�B�O�	�R���U�h�B�dl�Ȁ���ȁv���
Ռ�������r#�,���4��n�N��RpjN��Ȉ�8���\2�Zi��� e��� �\+j��#���/ndiy�������|�mu���mqQ(	����Y�w��P���3Nx�a@]QǀHq��>0�s���L3����L�h�
�k�N��\k�j'ra9lХ����RI��~��'����4=KK�SP�D����^S����R�����$
�i	�9lݽ{Ts��������%йccc�cc��Gj7'�;;͚�8g�m~�k�څn҃�ZG��h�Q}��Y� ��Z%�q���� �.�����2�:oXs��_o�5�zK5�"��*�~���h���t���037'fiY��V��K�� )f�Z��FB�ԫ녅}�5�1 ������h��z�]Z>?���"�ݪB�
j��9�v�N������8ۢD\LL�M�� ܋d��ҍ���3'$>��'ơe�����J��MVό˽{����8,8vdn�.,�� �F_��P��؊���yz<���2�*�y�ݙ4��E_[K��۹��(@�f����d$d�ͥg�&��h�h�V�?�o�o��yv�lC+� �&�&��� �`�ⶶ�M����O�0~H,�u�}�w�����2�3���NgR��]Y���bb��:��*�X�G�;��O��OKL��(�d|�4pQ�2��� 	�؜�r�t@jry-Da	(]�nAq�B#�� W����[PV�++�{k>&1��L�U6�cpr`��x�i��ʧ���]] ��T�Д��	��;;�;��[:W��z���q7�����9����~ke�mu�J��=u0�mheNʃ�8�Ϗ�Ӽ��;2")��C�Pf�d������|�T���h��f��b� �B�VQX�{���w���T9�7�-�tuuuvu=���*qi"c.=�Q�ǀ�|]4�g����Q�� ���=䀎�h�)09�bՁ����9klbb\�e@:W�KH����੡��C�es��C�k�Z'�gZ���t���s��B��p���@?ɼ��'�ɽ�����q����𓘀ܑ��s�^h�
e����[مa(F[[A��"J���;4v�1'�w�$����!GG�O2x<���4�C-�<Imz� �ݘ��|�G��*��S1��ś�Y���q�A6���o�x�-N�G ��?�З�k�EP�.��ۖ��o)�^��$���l� �V�{�n�gcc�{S*�4��(#Qv�̲��W�LZ�Db�X��]������|J�����L!u��Hčl7�Z�G蝨{��?�V��з}NXڭ�{��{�s.�~�n��˾a��K4�XZ\b!
��UH��T6���5�-����B-���Xg\+��t��Iw`�C�M�H�Cqw$Rsu�,e���V4�Ҷ~s
�^�h�ÐX�s"��$�`���|x��k{���6����J�����euf
�͙2�pɎ�!a; ���`� 8���&p\=(x�Epx���Gi
�;�z8^��������#����'ʱ�OojhpV����MgsvX� ��4�T�������4���H��-;&�� �)M:�����N��...���B��'+�А�=k�j)<��tD:q-���~��G�1 Zz��%�C����:�-���,�j����2$f_�9��cK{����Db��~���_�
3弤�K&����RR����M�g�fu��m��Ub������`e�`i�ɫ���}d���P3"�wD���ǩ}�Af�h�Ņ��&V�Q�o\Q_EOw (쑽�3,�������&��@q��ɚ��K��R/��~�n�����ď��snd��|t��J����H��iU�W�e�z��Gf�0����ҝ��֚�O
@�IQ�퀔k48#jn�<�!yv��3�c+�P
������$�&�5ɯI~M�k��C�Dn���I�?KM��ȉ�6����k�5����_����k�5����_����q �Cb�^��׶����_���xS/�S�v𮻫�R�/w|�Z*�,/-~=v��כ���|��|�h��w�K������/��r�s
���,Gp��_�9���{���>�o�7��~���:�;���޹��	~M�k�_�����ˣ�9�áwL���	f}�@ ����������(�Kٛ�~6��3��֪c0����� �^�Vh[��ZRw�}]��d�	�K�a�B �2�A���A���5�X��z�R�K�!}\��ϼ���6^_L]�pΩ)�M�a룷6�n�|H�
�Ļ�#{�m�Gi�̌},C���`���c�r}C#���?"w����aWO������$9i77���3��k9��f^NB�������"vUm��Tsr7�]ܐg��`.�G�w�6��}�I��.�n.�r	Ț����=���bp{/m cO�z�ԍ$�+�IO�
R}� �蓠o�q���¶L�L�eU���M��&�Vۆ��9oxZ����?��ق��Y�Z���cle��WD��a�8#d�S'l�����Ѣ�zD�rgXŪ��4*�R�m�WȈ��h#OI�]S�U4|��?�h�6�E��q�#Z<.W��FoϮ��Z/48U6��	BƙwLE �m�V�y�3,fz�Q���1�r�����&��޼u��aͬ.�����尡���~h�F���>�i{�;GmOGA �������k�_�4�����7��"]Y}[�',�]�P^V�u��I�M�?���E���4g;'�u�:�/�뒟��R�C:��x��劋w��PK   �|�X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   �l�X�4#�c  �  /   images/fa0dec76-8343-40ea-91a3-e67b9f04a458.png�y8�m><R����e(k��H��]I�+Jٷ,c箨Pcˮ�RH���RRb�$��3��X���f�~�������=ގ�>�{��u}��s��Lw�����-{�`0��gT�a0�Df����p�B���匱;�!���PR#x
.��8}�������%�+///��N��֗\��:��&M���`�c4T��{'�u��m3�,P&[���>������йt�����>���"p�Mʹ�������
�G;j�oz�+�D��6_YVop
k����Z�*�Y�S���=��~j�i܋�˫ɫ*\��.T.�*����]}�i��2&d�^��QCz���j���sZRR���ʏ��o�#I�R�C�k?�~���3����1�ː�@��M��P&y(y��}�5�t��s2X���5�Ӌ�R].ܗ��ˎ���3<��'0`D�/Y[T�4���T�-f�y���������'8�R�T(=�}Nsm�����<��]լ�!��/����&hSϫ�e�S�g�x/���$اM-)%�/&�}�����JL����xG�u��0�UvW����h&�JJg6	��C;d21�\Y��p=�^�\)?�b�S�x������:iE�=��II��ns�lZl�����`����o����=�z�����a��ѩZ��#Qr3��4�I�`V��߿���;��X�]����IRN^�7����]�њd��'����vG��|�^��i�E��b�����ǵ�8�j�&Lz~S�um���J!��&��d�C���a��JK?6Ycn)�3b*��~��V���Or���L��V2k1�n�g�u౑��5E�%d�Z�;5���k���Mnj[RC����=oH��}����tc_fآ-��"�I���("3�~�&�C*??�G��*gf	�vd���L��TVB*��9���̭A��?����p&yҭAѷ�:���k�� =sceq��)qX���ɴ���J`f����g�<���Yd�D��ϟ/��TE�%i:��+<8�� Q
d�ma8qln�XY��i^Icw�%��}�5��wu���^G�9��A�pZ �"d��k�c6��i��r�>�C�Ҟ��������+6��\�$e��;9�1�@�}���BM�p�����y�Eծ��QWGP`�����0;�K�U���>L\��32QI0�G�C�I@,����=��k�7���ONgA4�CX1=�s�w���r%y�g�o�:+�Q˽N�Dd֭!P�Ƨ�{��(��9>���C,xt�9�G�������(���E>�Ҫ8�uG��.G��_iƷ��ʌ��K���57��{qR�	#c�ʕ���2Ž�m�=���iZ��Bn��T�;��ƈI)�]�����Q2����ښfba1ߘ��O�q�(�f��i:�s���_���J�~=�@ eH-�f�Gbz���N�X&~��5D�o#b��R���N�Hfz���b�!��ZlO@�=�5�=�cL��a_[��<�f���Y��oX�<L5IU
�����z�q���Q)=��$cr�+++U��O��ۘ����w���e�[C�Cw*�ܤhņ��h���n/ձ��9������GM*�b-�/E�;�Y�"��8 H ��}"�ELκ�w�D���Ba(^/lC��2�fJ��6P�.���垑iڋ�����W��x'"�F %�H��Ųc�e��xX|�.2��!_Mc�!��@�3�&��^�|�Az�GGn��ap�݈�+�
�;�Y�bj����-
>"�J;�����7�1��KLT4�����s��K��o�ڍ���"�I��«�;Pt�{�yV��߃Ut�A-ODi~����Q��,sî\4ڎ�;��V��7���_�8K�\٧˰�
�@��ѵ��R��ا�����
��߃!0 "3G�:��K��&�Uu�PZ�%Iq=CP����I�5�Sҁ/�'Z
˯��������Wbp����-���� ��+P�|���Ӟ��vA)*��� �Hiru_c��9<dl�!�Z��0�D�=�(<X�ŭh9>��X7Ej���������Fb��B���9[�w7�{�W����Z��OM|A��!(gu�K{t9�E���r3�܅ jr=Z�e�G�
.h��z/��L;\���
я^�"Z(BE+�.%o9��1�����M��wO�T,;�ސ�g��|X^���ژ*_r�d6��	C�29(82��-Zd�M�6 �+U��p��{����HN�h���bEb�?�/Dl4��q�_GwD��Nlև'�a0}�6P�d�����~�h�˽���&��ʹ�Z�G�M�i(����<;�����FA�U�x��}�C�Co󎌅K��a3��<`�}����W���*��U�~<��'�;�P���=�ԠP��Q�e�#z�d�ovj�a�ԡ�%FFZ�'�j9�/l��9�'�I����֛i�M6>�N��SQ&7���4�K�zƁ>�K�����@i��xC,7�����>)5�^J{�G��nQ8������zJ�U�.EaQb�,��rkԝ������D�9�ݹs�i��u��8ݠL��x�n=A��Ä�m@JPo�T0y����z����ΑaRq=���i�3!�B���!��K}���"$��jb;�e�c�IcXRG=^)���²�U6�W���#F�c����SW����@����=rbݩ�>CǬƺ�+Zc�RJ���m�)n$,��׌��10Y�*}�u}B���dO�I+�oyի6��y�-�755=�dW!�Ʊ.�{�� 	��~���ְ��,��N!�y�L�i+�h�.��1���KƢY�]���� �1t���y���@�v�����W��د�v��l8�R4�Ogxv];��x�gW�14eu�Wi��9�1�� ���$Q�G�0�ԏ�V�� �9�����L2�;��v�M2,��?�}Pt�/�*ǭh
	��\��LG�tQW��{�ih����<;�|�f��~Bp��C���vҶz/$ c�w�������q�Nz9n�@����޵k�Ľ0WH�)��G&��Q!�ޫ�n�|�m׀P+�}�7��1��Q/v \4�?�'��N� �e�J@R~��&��EAG��t�Q���7�%�5~��O�n���hcu!���ޅ2!|���XX��jr�< �Qaڪ�3�V��B�7�8[�\؛�(����,0@e�!�j�1�� !��NK� v�T�w�JԬ���g)��H�B��3�&��(�7�m�u�͜������ �E��z�����͌����(H!JٞPq	h�יa��T׬����a5�V2�	W�Z�
X1;����rt]*�L�۬� �V��#@�gmd�	�(?:��N���}D����Q(��`�(���?���r��&�F��`o��a�쑾	����|ff���9n=}���B�?�"��Ȗ'1(�ozXw�,_$_/�������.�}�fϿq՛�ܻcK�}�rx	m��0ْ�]��gєE�z���\Ĳ��K�;u	$����ǴҶ<a��5Q� (l�+����uvzq7!:с��6v�C�hQ���Yyjf�ŒڗhNM{�uKhiiE�Ɋ��Ud���!�$O�[��r��P@h��Cssx�3�=���VvWk(�[Б�hF�\!�{aݧ�R]Sf$v�Z��=��
���ǭ�0u�6��L�@��A_� �3��ߊ���O	��fSH���4%��	�N�yۣαg'*	���kw�Z����t u�B��ȸs� m��:]�~���)����3��p�Ŝ6s�BÞVh�<(S�o`��5��2*�4�E��Y�?㊊�n���Y[[��To����¸ �D�����}��a�\�O�{)�R�%"��p�6�y�G�=���F��S���yȦ8�N7Q^�#���ڂ��,О a FA�ݯ���M?�R"���]��F�žP1��&����k���X)�9b"t�(�#�F�Y���q�+q�����a��i�A���1�,`�/�y�W�l
`ة��f`�����U&nﾯ�_.���f����4Ћہ�1���T�_��W��ܭ����c��E��1�TW���x�@�b���(�CZ'���<<<l��i�G|t������EY���:Ob�ģ֙�y�f���r���taz��6= ��"�"ܺ N�H+��$��ׄ'��'�n��������bm�A��G*��`ǯ���.8V��	���pɜ��6d��uY���2��� �`�V	��ѮW7��	���Pg�|�oѦ��h�]O8)��i����ć�@t+�3S?1�7"���zY��P��3��r����g}F�[��@�3�AL�m#�Ͻ��rL�Ac���ð�V���=��E �Z�Aqi27~7C^��Ѿ �9q�pK��y5'1��a��<z��W&�w��7���P�	�Z�n:l�5���T������tbX�#D Ii���v��@�P|��uVhc�m�lre�_?��?������^s�k~B����f�C��TB�a�� 0Y�A���r��&�Ò�`���M��P��`B�iHY>H��P[h+�z�""���/Q5��R�@���������� �ϣ��J��`J����\՚\D��a���k�Չ���-��e^��n*z3�=LJr�H�X�Y]�]텊.OыZ����Y�a�P�=(��Pq��jIԛ���	�c�F�.��䈯��X�od�h���RC�C��Ϡ*���D�H�247�8������s���/��5���aT����yo�?h���1�Ov(|�H���`����#ی��G��~�ST��#�/ ���h��.�h����� �y� +�z,��:՜�ԥ������s����� 8��������O�{e!��݊����Xg�䏰��h�=0�E`wU�h�̖��V.C�;��aa��--ϔ#H���h�
;�-l�QiC0�y���p��@6��K��T���|D<����}P��a?MѮ�Q��tu%���L�\]^�`���ct%�3 �C;ֹ��	�Y
P�9���P&��~�Y���}@��"IC�V����1z~~�����?y�(U���ͣ L�-�щ��e���0�@�TW%���9D�)(X�m '�h�xH@�������)3��?����K�����`z�T��� ���ЊG�t��L�Q
��[��[:P�@�z�=4��Un�*��af�f5&.�89���Ȥ"P^��f�]�_�7�y#�.q��ioz�3���Z�*ݭ55b���r�wѣۉ� r>��S�G���P�/G��N>jU��8J{:](����jRU@�iO);XPU=���t(�T� �8d�k��K6����Jf�}4��Ti9@��(%�q  �v��$�C�O����Q�]CXɑ�ri��ACvW-4��L�y�i�7Ȃi��U��u��l��Z��2��*p�&KeY"]GP(���
�VV�4�'��m]D��`d�c�������Y>��>���(B����D�݌��Q�0�ӌMLd� �����V
U�V��#i�vt��!��� *'�h	ڠ�.Zh��?�ߪ�=�p�L�wX�.x�\�p����� '\�����Q47!V���j?�a�2KD�t	A�T���2M)�J� �v/�o��E�c&�ke���D6A�����e ڲ��n�@Y����A)�0\4@�s�(2}#�
�G`�SQ�o��K�/l�$FgG{3���?�>�����0y��#��M���7u6���& +��(� ?��?�
�tQ񯾪�O��W_)o�?J�W,�w���+�������AJ��W_��(���6B�*Ee��W,�3�i��(����������������h���o}U,8(u��+ڑ����R�}����������X"���9�'U�(�7ا��-0�*P�%��H+Zbd0��0S��"��T֟�>�V`����b��6�>i��u�fs�$�C4�h�PF�#G���D��B�nA��Ǻ�R���5潴�*�Ǩ�R�'~B�t�ϙ�Q{T&�t�TF�)��9�ʂGN�����kH�O����U�U�y��.,�/�)�;:�Q�L�0q�I�!~`jbb"&�.}=r�(�,h�tuzK!�V+U�T���Cԓ��z��E��ˎ��FV;�dAH�z�?K�jeF|� N��R�����@�5Q^8�"��82�-�D��m����IE��<��k8]��/1	Ef35$K�۪֣}�c��[���1O��m���8�`rs��k��A���+��҅^Z�n�����|=\R^.w�~@ͦ_�_�ꓡ���Y����o�ǻ/X��>��(5������4�d8A���ӓ���+S:��j��~����5��n��9�Q�{��T��l�Q�v}���e�'x``6 3���5(zu���� 1�	���S�}G ���9�[8�*�`�n�zv�LuZ8	Fi"�GP>dK���n�>z8���g��(
�@��&b�͊]Z�ԾE^d�����g�F�#VI�Py�m h����-y���NmA>���	��#h�xHw^)�؝&��e
�yHO�����G�9]WC�.����{�$M��U=��*
u����������h�hTT���|�f�4��TOF6�2i>�K`� �t��Ga�V��;}.���^�1��l�tR�1��� �Y����t� ǤD\=������S\���;��e324��`4:T�0�N�Lc��?��_X�ۇN���\����x�S�V�]t�?��.\�\SC����M=,�IG��|�=9��A����"t���O�vs/-BDL<h���ϟ?���JP#fh�i�q�S}�N.�޸� &�d}�����[��۟#�<�-���7 �ѧc9:����gRT���a"���7�֪���8��eB;�d�H�}�@��b�]YNߐ�"���e6���K^�����#,Kס�9�o�Ţ��t�!{�`�$R���?ծ�D�N4�J���L����i"U�.�E�$���R�1��=CN���OWW/Qn�6"]yOB���S"���T�f��a�����XW�Iͱm�X�v�67{�&���]�~���ƹ�P�� �C����t{38�0�IB|����x��g��F�Z�Ph��Aߓ�4�Tf��h�E�f ��i3�	4U���qE� b��/i?���ء:ɠ}���P�,QG�Y(A�.��A�V`� �/���$����!���1���C#A\�����Ѩ�uX+th�A�?��)q?�.Zi�@k?���J1�� �EG��%ʳD�����c
��V�h��#���@>=����V����� ��"ۋ��Ѷ�*��hL١,Z�����Eņ��pF��^��6:���Rd��v���<�� �m}E�3��:�B����_Y}9u����#-]����PqOi�\OTK7(˦�eS:& �O����\������3: ���R�yiG�A�@��/��j��p���e�)��� Vt}��M�* ��S ���J+��)���	�UFһ)1�Z�@�5�t:��48w�?���.4�V��6�?밴��/++��J��ӛ!T׈d0F�O��/ϛ����2m�����8�&(�i<�;������5j���6:��l���E{���GN�rٕ���i���Y6F�~��~������CXV2��tD�F���?c�j��_�u����XA$z��K`YmA��_����q��d#��Y�q���A������t�p0��z�"�֣hn1�ڌ�X���Sy�K�e����~��1@��~�ut�&�=�w�OF��ܐ꣈~l�}�N�ڰz�\�f�"�!0�#0VI��f4�����hO��O��:y�s#���#K�^.T���@�) ~�VCSv�	`�:�� �(�����`^X-A�b�Ġ��������3dAU��������P�!MQ��ePB��ĳbe�7���/Ϊ� F�ѳ?����UA��yTX��c,h'!ڗפ����3��7�������eXH�խH� U3:�z">�ێF����ޅfCo3b�E+0'���PT�cz��iJ6�Ԝ3�)i��f�g&A��AߙWﺗ1�iI��{̼����V��P�KF�	j�!b�6����3Bx0��&�j�!0@�0�������^R�"�¯��6��t/pL��'1����~&�I����/���53��bn�e�ا�Aw`0Ok�H���+��E���m�Uc���]�z�%�%��5s��\��b�6b�<�t��\�<3�4'�ڑw�?nx�?��<3l��}��0��~�\��[�K|�k l�(l��0�����Ԇ�T��5��5e^��������:+���a�a�#h��**d�����W��������@���L�8���x���_�O�w���X)���I)�Imkw��� ��<��W���Y���`�S�I�z�	���L_vg��,�����
{�=նv>���llԞ�_��+�����%����ϑ���TW�=L��䄵�l"��Z��|�.�������g����v�g{��U%U?o��%���J��e|���}��԰�>���\N����t�j7���=�\�!H���(�KP}�8|
ԃ�[�����I>����+�'Nn�`��m"�Pü�Uy�	���!/@��6�_�5�ɮh���$o�/��rHI���?V��?����_K
���1�Ad0�B��9���&>�Kz�/�j�3o�����V�V=T��j��q�AJ�7�׭��p�+��j�������2	7�4�/�����rO�8����u��b�e|��a:�B��aaR��z%�u�Ej��l�Q?C�#��]o�^pHS
̅��g�;|O�V;П4�ϟI��f/��OT�R}<��f�:Ȣ5\ xt��<A��^������6���!<aal��!r?6��)��'��3���46z�s�[���4K[�[T:vD*U9��-뫮����T<�{ږ��Q��;aQ�5l4g�G��ң��G��KP�Ҽ�%�m���31�
�-	�vU]1!/d�e��[�� �b������K��w��;e��JfS����^�35�bDز&��7�U���#&���(o��jym�ʫO����7��m�5��(�f�k����!�2}���a��h/��M\�����ٵ�3���v5��^��
���b������1�
G���u���
�q������"Þ����9�a�2<�����TmՕY�T�*������1�g��jԭO���F����r�,��������y@�C�\���X�VO',����]=W9a�G=%��	�`ˣ;����a��8Տ
;��Ȩ�}����������S�ől�Ƹ
BX/��;#-!ԯM*pc�E~�� 9�x�bD�m�G���9�⸿K�wF�gyW��82��-��b���%1ZQ�Ȉ��N-ڍ��K)��8Y��[a޼�Nb��!bK��W��Xj�NY���ğ���V<�����k���Wی{oS�l�^�k���`�Ȱ�z��'���O|�\6�Egm�M<w-�?�7�����	�q�w�u���V�Ġ���0;8��GL��rЊs���n6/xo�{����������F��'mK�Ƴ�U�m��m�Y!	G���
�d�gm%|Qf(�W�;ȁq�e���.��ˎ~q�Y�=J�מ1�T�?�5��I�	���Ab����p����(ki�F����v�9i[��<?S��A���Y�{ʊąQ��� <�#����e1�dGM�6zLg&)3Ti/Vڍ�Ma��h��[d^�f˄A�L�sU��G���[u��6[/W�.=��g_�����Yڀ	����^�;\�LV<�]�1�:���yN��S��7�MZb�=M�<��|(��B�O䧜��Ģ�<B/��\�Y�|?X�OyФ�%:lc^�^�h:p1�;���Z܎���$j(�ˬ�z%^��//�@�'��uUK����Y
Q"��\��e���#m�4�8���%���OB�T�Q���B�m^܂��?�� 	P�͊�6Y^���P�`�T^����7�x홭4[bNlڰ���D�F��5��ۘr�~04S���R+��%��.S�WR�<�� @���*�g���V�S��EK(��񨚿���II�f���d�6��MU�ub����K4Qc=50`^r26�YzUo)�E8!�#L���eU�[�ŧ�Ү�����6�=6�y=8ÿVNF���r�^*�U9�?%_#�	���9e��ep�L���n�*Fb��N����'����� %��G�6�;��X�r5f�4*3h�X�C��4, ǌ�|���Sʁ�xKalH�L��5���S�k)���>�+���*}�&'�YoFl�����}k��AZ����l'�3��w��D����,/�C�i��ʐ�ly�2^OH�nI�aCB�x��>��2~��ժb0{��j?'�[��9�蕑�'�I�����{�],o}�ś]@��m�0����k�9�/���ǧe�U�u�m~z���)EM�v�L�Pe5.��նIA
	]M�l�����0}�G�j�����2�"�~�"���|�D�0��å�~�*~R9k2��/���CN}�<}��퇇�ɳ���hK_i�Yʇ�:�^��2[���O��>G=Xǘ	�����h��T��dy�_C��,a��lW�V?�_e��{M���X���^%���Z�c;� �nI�)=�ҥ�9ӟX��T�/^��q!(��WAfbW��?b��_yfU�(�7S�_��ܐ/�p�8�g�ra��wm���H��
�F`��S9�|z�Vym�ߖ<��r��2�t`�D�LM@?���O��V�y�p[o�(����|�n�^�$͡�a�!a���L�p���:'�Z��Ǒ�$��8(5���=�<��L'wa0.=�4հ�G��P��*~4��6_���u�������Lwr��ϟ��i�?�Tf��ío�V>7�KJ��K��/;mSn��n�H&���wM�ײv��ϻg6��X��������4����S��֦���R�5N���A���G����F�P�5���b[���˧�.~h��}Lͥ+U�7�ٳg�xR}�ШlJ��n���(�1k���]>���W���VNW:_#����J�����ŧ�ye�mf�:��W��T��L�ּ�2~�LJ�_�e e�WϽ�Ro�L+,�Iک|�|J��Ŷ]��~}�(R��z���Q{�s�!��e�����"{�ӽަ�L�9�VCC���7#=8Rf�g�\����ֽ'O�TŘ��5*gȖ�<W�SL��dz�`0�b���>?��ZQ�.'g��*�|k��g��Q�E/ε�W´IO��焵|������9���:W�W�����0�n����r,�J�R���y.���O���w��x��r�����m���V����������M](�06�(��$&�cc�abU��騼wg*lC��I1lƤ��V���mm���|�g��F��l*{�m�}٬�rr�d�$i�>�ڃ�\|��,i������*����<K��.ڀ�شN˵ӱd��vl��Y���<F����|U5��A#0@QT�`�)�7upr�w����A�b�n��0���e�Ƽ��r���'b����3��?vX�CŞ�?�SLk,��Zr�.��1��|�K.&6��H��f-�D>���Q�+�zx���].�z���g��7Sg w�D\A�������X�r>�5��Whך��_�m��}�ر��?��{��Է�z��E��ZB�!�U?��~�%N�ZZΓ�T~����q�^?wpGfR��w��W�0���;Qg�0��tl���lccg/u��&h�h�@+�R��<ϟ�9-g������I�W���V�<'{R:��*<�=��I�Z[X�	���f?���Qd?��VY��j()!�n�[�V-��g"�zv	�<؄�'lߚ�ej�4g8*X�1K*(L$��|aZ"�0�4��ƾY����wa�|�F��ݶ�ge:���ٴ���X�0
b��HJ#�r�����55]yNS��C��66�G����/���ڑkh���I"�����n�U��Ԗʊ�������1�xL����+gb��1�c��cWľꭑ�lGR|�[��4�2;K�Ű�A/�&{~�.Q��|l_�74��)�p��$�Sd)�C���>)��jVy�|C�I�[�*r1g7�	ě��gO�^���oN݀ѹ�}xD�G~�s�Qz�P�iSգ�o���2f[ڹ^w$�ԩn J�Bf����˩�Q��Y0\&���"�GGf�%�f_w�,'����mX��X~�����M����4�Xn���a��K����L���3E�M�S;{uf�_�	37w]��v2v��d��H%Ӛܝ�����ܫ;���Tuˈ��]�e��5mw�<�a�����zK�d�G����82,c��f�Z]�O���T��5��u�g�C�9h����H%��e����Pu�5�t_�yܷ09��(T�O�ݔ\E$!)i(�Q���V)��J�Lk�;���㻚��QKo��ׯ_-��㯐�?�a���>��h�y�����_v�w2���LkGL���!�J��<l���({50���5|�����
V�Ja``��|S��uQQQ�l"�k�����,����fu���qo&j̘_��P4W^�ϸ�>���w���6�'P9_�?�W6qm7��mf^���lP_"a�Ou�t�؈��l�����r_����rb�@�!cХ�;F�ύ�E����B�ڊ���`��b�F@~��)�����MǮ�w:��D�͜������x�j�$�/�eo�^{��hr�Nr�v�������6P"�ք�د?rM�o������MθHe�V׆�DI�W�?ީ��f��e4i9B��63��v�iy~\�m�J��x��T�;��ǿ� pIj&=pOe��ůR��V�J�?)?}m�_��&��J�e��)�Qk��L�r�='JW�NVȨ�:�p��_	��8<u��y�nty��3�oIR�����O	���(�DK�B��3d���S�J�}��6J�K�V��_b_��vt��B7�M��?Q�Ѓl.e+?
`"aϱƥ�8(�m|�D�,=��ՖuP�|���Nm֭����Ί��-��5.Ĳ�n%��?K���_�>� �2�mQ��Hj�z�ོg�A�Yϲ��T�An2G�H�8��͕��~�u�Y��_�h7Ai��p�=
�Z)t���d>��9��*)��1 $�koS���|➛>�f%9}1ГG�T��y"���]�<��m��2&�d�H��p��k�S��VsM�j�s�z��o�.�	F̞K�%}(_-��#�I� ������`����m+o��b`3�fq.�D0+�w�*O��E>�+���}��s�#�W�XԤ��3~�V��3x�Dޤ�,i���M{O8<g;��&�]R��:"?�${��&u<�3�����﷿�-~�q���HIo�/�=a4�7-�<�_bC�mO�-�|�7"ul��fG�UG-�p ���1���W�2`��D�+�~���4�0��3�W�w����e|uI�-�XT���܋���T���<%�������xr��ܨt{
����ƅ�-.��v �D�<��Y��&��\�hC�Y�3;�J�X���d߉7P(�7D��ne�ՙ���K����;\(Tֶ�ʢb�ʴ��6tW�����r��������KEIy�y	?��~�^�!��G�Yn���bn�
D�J]]v�5&��<?����@����zۊm)<��P���ה߃a��3Է!� ��}usm��P3F�sF��Z���mGN��Β����ͳ6�q�ҟ�M\�Պ�{��uoQ���`����P6��˓UU�.��8��p��iY��c��Q�
��rIIr����~/z���������UK:��*.��H�&���Z��̓

L�pR�L%|����	?I7��ZN��k/�^I�6C��Pa��8R'�F��b��S!�1��i���E6��K҈k�3��#��� �$4z�|�sz��QU��DY�ǽ��O�uN]z�=C�J�f�>V�}����8�����x� a���G7��..z����+h�Lx�_)������}���vU�!
�Q�g��������`�7�ϧ��]k�>c�P/`���2�Z�WL�:L�{��� �10 �^_�=e�%�V��5c}o~��]�����$�ؘ�.��P8t��Z�Ng���ڍ�U�	�&�7��=���a�	&��ԩ�ן�:���oy�zh\�@��1#�V;O��no��ɱauG�p]m!�bu��7>���z��_nZ�F��D"�~�|���d�A�q��}C�wo?���*]6��b3J����in�G�w���(I�.qn% ���Ǟ:���Kvv9?����Fk�3�=w�ֆ���_�3�=ހ�`�g'L�)�P?�r0#���Ro!y�M��ݪ)�����=�ћ).�^��]q�8Z���<���҇[��&�+�Q�m���5�9�b�Ll̼���5#C^�Ey.U'θɷ8A�.��Y����6_� 3ՌlP]Z]�	*S1};:�Nv�;׎�8�$�.������m/�c��4g������sr�V�-�SO�7�V�b�����ܾ�挍��Z��gh�<G�= �[ z�%���V}nIOb-��O0Za�T�}��}��ٙ�*9�T��$����l�扯S��x���l��Px0ȹ���p�?���B>���!�]b��' Dܲ�j���Y��zs�FOo�h�~�.�8)p�t���>H�((�/=<5ݢ�`!RPS� ~�ᓅB@�L��_���B�f��+Ѥ{t��KC�,�#je}!̯ps���=U�#�<N_��w%X���,ds��D3v^�#�s\���+lu�	,�	m����ǯ�4ǐe��b�5�?T<mG��<^ՠ�F[=|�mfZp��}\�����N��C{����ͅ���z~u|c����8�+6���Ŏ�h�x��)t�v�+�����M�x��ty�����'^!�-,�-�c��+����_�I�и���hE�F������YS�ٲ��\M���{*��u�����+��$�J1���'�{�P�a����,��3yO��3e$�Z�R�и��݄�'�'��R�ڳ���8�W��h��o�{b���&���߆��>���e����::W�Y]۸�b2����܋�M:*ܜh����8�݈�f�N$��Te6��RO������wSy�@a�{��!��z7F��Ǌ��@�2^�������Y��,��1!J(��#��a��������)��6�,t� ��o���4�l�{�����5�Aƭj��Rԭa_�Eb���1��Y�3e=�B�6�jNfˆ����5�����n��W�#��"�J�˛�|�%!����@P�bO��tΩk��33�����A������$��4E/�3�ZjMU�W�A~��F"�#���-��:s�>?Z���wk�^�,���<� �j/����]�47�U�u"J2�'���=��ѳ����!��'�Ж�k�G�W:z�a�5�2"�@���O�bC�-W�9g���|3�S�;Iӌ�/�Q�PyrhC7����n�+����I~��fn�j���8��~x������c���k�;AoDQ�8���Ġ���S�DdF�7�7s?@l\�Y��+��2(��u�6[��O�����d��Cnο�����$��^�d��v��*� ��Orz��"='���5��hK��]�zА-�3�bH>�C,�dė�	�mx���S.-!��bK��yFg��jWܲ�]����|��䙙7Mʷ>�E���&+�`���m�Ɩۀ�����;��������D4 zӱ�G�mN�����6��L�O��HS����so&ގ��HB��wr�S���ԟ���g��")����Y��z���}&� q���\^�ry&��->k��c��Q�'�Ɩ���8l�kZ��L����4�|~1[>t^�r>�M<N������y�ac1�F���GM�ß�:��	S0�+�'hE�'Q\5��=ږ���s����s�K�`n��%�UƯRǎ=ͯB�mu������H�ї;ȿ��@
||0Z��aT�؀�.�EmÀ��w�!�7SáG+"�G� ���1���AH��O��� ��%�c���ey
ax8)��v�?�3��q��Z%��-��9ȧL`�b~Ň�.���v~~rhä�v]�՘�gD+��؟�m�+�Qq �"�"�/И�|�w��h��Zp~�����N4%���+�K���簸G��!y�St�H�٩u��CG�p�۶c��>���eh���,��S����W���I�ig�Ų�o��ȓ[z:e\i�\!�G�}	�^ؙGr�u5'�m�` ���Eڙ����N����H���W����=��k>��}��;M ��yb�UN��Y���@@�}�r�3? zϿ��qӮ�:��;ώV� g+��<����a:����1U�)+���	��ht ��<�����aki�s��fX������D��*qp S��7�6����}�]��RWk�]����H�� x������<yV�Y��/!-Ws&�X��C����\����( VR�H�`�N%�(�%��˟%0��	I�W��j(ɜ� ���9�.N�ΐ�l�'�h����GX��"f�4��G*v0W#��ɓ����/F�0�E\>l��#6�l�4�o��B,�6>�k�r}A����w��9��������I�-��냸�%��E7��+�]n���]�a���S2C[��;����=�8�_w�x����+���x9�\����x����A^��el�t��.2�o�^��y�3�`�;D�߸����c�7��?���ya��˒�ի�	ㆆ�8@��w�5���<���sҿ,Ϙv���.}J$.�Ҝ��V�xh��_��_�q�B� ����j��-ʤ��o�$z��U��/m���B����t�.�{�m��FE�v��9C���� ����222��<I\>�_]�����4joŽ[�\����o�7�"=hmm�i-�-�N缡a[�)y�]XAM9�qxw�����ŝNG�9�� �#��+o�+����:������'��:��ʨ��,��w~��T���DI����L��}�aGN)+ޜ�w�7�9#�����̤Y{-��R���[[�tf�\�{������ʔ���+6iu�h��)E�?��F�ω.R(7�x,��YU�x� �y�6�/K;U����.dZ�����i�L����^{�x�n��4ě7R7oX�B?r�88h��f8a�^����E�L��疫���[<���b��\�M��5���T���J��'��ԃe#��2]�a�o@�d�mB,���V`r�d]���OC�؆g����zT��B�<���B7 �0��m")n��� <ŗ�3���1���2N������Ջh��`�G���R�k��G���¼���ޥٟ኏����^�3���W�] �!0Qʔ��o���������=~���N�ƶ����įG��=hԌ)gk��RZ7d9��̋V���T����&�:7b���yI�3���t;����e��7S��}c�N9��x��f�k`�+�ʚ� Q�e݂P���gW@��u���ю�.�#�n�?����|J��;��|fF���n?���YdoTI��E�#z#|�1[��l�p����&͛0bi��G�xv�g��9��R�]��5�Y����;��=^�X�?&3-��<䳿no���a7C��V^�u$�kJ�I`ِ����E��u�qF�_��@HH_\�`�w�>ba�M�� bh��ߝYA��+fh<<Ģ��H�Nr���l��o�T�����;�V�/Ϗ#�a��w����{�B�!�1_��x��̀�4)e�N��q7o��Aڴ㨼|JB�f���A��p?K��PϏ�1�W��/�~�tU��[hSm==Z�o���$h�>SNLM��Ø�!�iͲ����w�NV����e�{������7|6ָ)�'��6 '��8����n��F#)�Wi��\�埜��Y���+JK�*n����uߘ���z��u9-S6�4IYnd>���~E#�ygLԙ���W,���T`�|ײ\jza�������?p�7%���=f�mso9�񣠠�[�����sh,��;��Ȍo1i޵R������P�m���
��+���I�Yי�"�5mx&x����¸~Q?�e7�W���w�v�ZɨY�2Ly�(6�l�a���V'�g��l�ҽ{���yj#)�TUY,]�}��>a9�����9�W�غ<�u�O�]�� pd�A��,�V	ϲ�ޤ�x��i�J��J�ulP���Ƞ2h���"a[�`��0O��2�	�۠��D��ѣ�"c�i�P�$�B !$yu�@��o�����}k��CU��w���v�s����3f?�N}@6�ܟ�`ܤ,�%���n�L�$�%������)<�v���*QAS���qf�����gU,o5��9��<�+�F/��}[t�������
����v�M[_�x_#��(ѽ�NY��q�J�r:�u-�UW�����}�oW��U�0'�5S����t��'vj� ?�����g�@G ���'#��v�c+I��4�Aǰ��ǎ�NG��NYN�,�Q�?&"�ٱ��"�}4a�c=S
'��1uߖN���k�}��I��7�P-�sT�(j ��q8�U��2I�⅌shm��ɼ	��r�#m1�Xli��$ߤ�@}:V�֏����M8�g�ɓ'���8P��(��rJ/4����+4�'�)��떙Y��_�pVDA� S���me=�w���z^(�� 0q4:��G��j ��h�4`/����2��3�y��)'�N�p�8o��YS��X�P͝�o�
�@6��f�&��E4An	����c���Cq�u+�WѲ��(P��T����d���%�f>���ֲ?p�f�B%.Ge�����~�~IB��%Mx-���\��v���F[^�xI���;��#��Y��^ps�|��C���7m,u_�� m_���Q���ތ�k�~������Ԩ�'݀�Foet��q8)�Ԭ޷&?@�<J�@!	�����Zf���:�`��ͦ����s��*M�,eЯ��{�&7�8!nA�S����˅u�+��4a�Y���F�H[9�����pzd�{��R2 -`��m��EdJh�IL�ګ�+��fO�g�OE7O����B�p2zp��V%�����U)�ټ���w0����q�H[-��m���)5��C}w��e��}3g_��b~t	�4�m�; 6�/�ub�H�M�M#�s��e�ߗ�����9��>O�f�By{m�~e9"��t�����?nh�V�n���vպ�g��͑����x�6.�H5js��3�r����A���Z-�uV{@L���Q��:5���ie0p��C��~�O� 4�d�Vp*=M��*�����B^���ޟJ�C�3��*���G� =��F��uj�F��wR�B��1�£�hn�=p��8Q'��?��Uz��c�w�Zs:.��?�&P��O6��`���6􁙲M��HԐj�ꛛ���VN�V?@}�K�u�.��9�A�>�%b�B�iD�+���� ��d�W��v����?qV��Z�7���' �I>j�{���2|@s�K�m��(sږ��1Xr�}����S�����4��s�,��V�\�=`�l��^�E�rʀL=����M>�0�������5�<X���2
�{VS���3O5zi����i����3���5� ^#yĥi!��}��\���ō�F����8�۸`�t��C��Ұ�V��  ܟ �쟇�ֹ�?�p�&*E�7�W��j�\R��]`j���mS�`�Ch <�o��V��ᔿ��4�Cƭ�e�@�2����)��6/�,��������˺��33�����T�7��<M���9L"��x}�0�h��Vc;Ӧ�<kq]�ǜV����3v�ݵ�m�p\�U�G�4�.W���xf=�����"�P}���(P�^��N6A�ڜ�3	��q�1M��h����<��F�+A����,�N�T�|̆vnh��$�:���������^�/������Q)�^B���6`�p��99��'��瞭T�wiM��n��ar51ѽ
l�_]ߧN����z�=�&9��,���MI���{��K�*|�˝����И�D��B�ځ�=J�s��4��<��LRB`��@d���}�� sAR]�)�`ߪ}`�+8#��`M(lZEͳS�f��j�3�@9��No�ny�`�wx�0T��S��!5Ģ�~����zC�.�A��j�O�6߼�l�I���$����y�>���Qԣ35�c0P�l����\ܾ�B�.���|�=@��E����r �0m�Q��'N��k�ԫ����f|���q�1�r9y�;9B���<┩+KV��Ǵ�l��K�=|.Z��]�[TTT��%i6�N	�AgG�oV�����|۱��d��V��b�H2?n�µ���/=ud���Ө.�db��>is��h=�&�<�ت��!?�m��"~�x�YYG铚Y֠i�$�X$g��׷�O��t���IM���rGS��IH�Yj�g��5�P�%�
�碣���w��l!���9aU��+#�Ԧ_�n$�����$���{�J�U��|��m!��|��\��j�&�F���c��R�Ŗ��f���l�]�P>�h���~+|^�p��V㊯[��k���T��t8���;�}Y��`�L����"������y���T���$pn˩O��n\�����V����M�Q��g�'��,���̩p����.یTy'Ī�i�A��F�:�#^�\����޳j�Bѯ�X��&��sJ[�\,����pp7��� +cPt���2Tc���Z�7Mcڂ�ҮR��6sT�Wr�OJ�0�럑�R�թɛE��p���G�e�,�b2��L��ڲ���V>�������e=e2u��9
_��%�}�}��0��������^X��\�]£��$���:�N/2~�L�H�V��
�D��?���G�{�DU�����Q#�*��G6	���ك�f��'T/}�Q��H6�MDLp+	��s��nH}"���2�Y���ٍAߤ�8-�}���2��?06�=K���zz���H�dR����UږpꈗJ��.�a�A����W2��%l=J��i�����^t�?�.�m(����F"������ӘNQ����Db��J��	e0$�ë<t��'�	��L���������	�׀H�ˑ�|��{(6wdK}"d��8�.z�&/�
�y��f� �_���7_��U�-d���o��yz��v�G���F}��t��t���� s��宴�Ԩ�i�UwC�.ډwo���@��^|�i�{�B��D�$ҽ��|��2=ֵA��81+ܱ��݀ �N&���C�6l�'�Yt h���py��,~(�F��k����a��	����rb���_3.�<>��y	����-	/5����SM��V:?�e�;n(���Ҁď��NIW�$���܈�ML��L��]�^zbs�}1.�B�[����6o�<�-���2��21��U��@E%G���"Re-E������`��wv����L�*1P��sa��$,\W���d&\�6$4�elr�C�F�rA�M�=�C�C�+� (�*�$S�b;�і��,oGH�x?)��l��Zܠc|/�:�g��_p���|A���1�ҥKGI5���򂍐��_>� ����(4��G9rF��@�1����S-z�G��el���D��-О���Sk�;�M��Ӣ�a�R�Μ9#
.h�f�'�n�%VY��Q�����ZNěׯy<ºE�`�r��Or-)z��=&���:%%��FG��8/&6�g��A��=�1���+�;C��)m��k�~� r��=l��nj�*((I2}���M !o�H�ݳbn���܂^���� �+�`=H��ئ�k�/vE#Z[��B�1v1�\���ŷ ��s�ơ�Nۓn��Da�N}���o�Y[�͂v<x/���3���>�1���&0�aqd#��(��bI&v�3���&d�w���^���*a�C>���hv��	AyHe!-�9�)n7�������'7�jb%`�+4�t��s*0YM[11�ԡ�E�Ba��+���_�Ro���}�I�Ii��%�j���'p�Y�$�W�;��6E� �tH���E�e��`�Nsj��AX� Ӣ�i*F�i�������e�u���A��X/߆��Q�`ы��x�IМ�.Y�d_�reG�&�,{�k;fJQ�f� ���%�Ѻq��*�^1M�y?6�v,|��"} n��T��|�|sQ�v���H@ϖ.�s��X%մ�a��!�p��ٮY^��-)=g�*@)��e��X�����#e�J�N�"1I��4u6rpVN�hp殌��ջ����ؖc���R�{��~?���c��'G}8�A3��kCYZH�����@��.�^#�9�Sqe
��ĨV����MXs�C�k��y�X���vz�)mQ:�����y�����J�_��p�R�7��Y���X�7ڣ3S��J�]�Ҫ��~�x�F���n 
^D�R��e}ϊ�;j�/�ǾH���;�7�'�5��Z�k�3WI?��Yq�;�s�o]��Z�l��!�����hAkL��y�#Ī�6��ۮ0�;��Nj��EW=�#�r��ן��`�mjF��p*����o����4��O�i>��ђO���x���O�O�����eh؜Ȫ��ut��1;W��l�o:s���+���S)�E�2���ix8�J�0���㦢i�n���yf��R���xE���fRkA�7�"A�p;�1��G����u���T��L����~}.#	�~8�Wj��~=��=kK2�#�x���F8+
3�|�J��c}�YwKKK;AS7�Ė�����W�?�<Z�.��V�N��SG~��������#�vj�e��,=����R��e��n��G����g[�].~SDz���܂��d~�!��yWWW24�TV �/�kS&>"dPZ�������ݟ�=��Rt��G�2Yw��:X����p�%V�t�j�E��'�*�.��d	��!�����T�sW����k�izc�eb���Sb��Mb�
���WL�4����&ȩ�G8�q�s@�໇G<bų���_��p�rym.)��.ssɵ��*c^�Wp;ɁQ\:���_qL�z��s��,������,U��8���@�W`NvS��Ȑ�5�c�C�>�?�%�*55�l'���	�ik���r��1�������]�����X6*�aI臁����r�u�d~��0dz֋���O�L��67$/'7���*��G&�P!���)|Q݋/4�%-�0,��״ˊ>�=E�g�"�ܩB�(�,��ov�����v��	���TU�ӧM�y��/��s��F�������I����푲��B�	�!�n�<�L����&N�<��r���ϸ�Y$P��y�]�T/>�q�'�QZ��~5@�O�r�|}�X��>rK�$��cO��}���r��F|~P���EY?�Aj_Լ�ϊv��k���� 1&/��	�0�ƘrA���Y�H�U���S\/ d�4�7n�o�<FM>������W*w���ޝ2�g�
��	6좔�y��S�D�Uf��s���6>>.1%/������Ç�+3����<���6 �Y��o1�J_�zU��4�a�<e�DlYΫ�C� <���g≂��~�U��8�3V���)qi��;�D}V:�C�Mj�_Fw);�Ҥ��X���1q�G������^��{8��< n��bL�o!���:�W��2����=+���f!��i���Q���!_����]����H��IB�8�1E�֕�]�y�M�a2~ոH�-w��u�I���g  ��7����gf�R�����:/䕦 O�sjO�&>�P"�4=�`�S̋
�^j��`^}�/�$i��ך�kcc�p�v��5�h,��v�+sh�Kd����x �)�9����b�����,i��%4 �D=Ax ���߿Z['-��� ��Џ�"���L��j]�+ˈ�X��> �	����Ў1z6@X �9&��z=��c�G���4���S�,�קԎ�T�i�}L|A_�V�DEM/8��nIh��7�!l�|$A�T��W�զ�+�&���}e�;q�L��M��-�I�>�A�/�~��$���V�-Mň��r��J�j�����t[Y����0@;�e�}����@JW�׿�<�e	�v�x;�� �xjqh�3@�$ �m�و��Y�#�HشPS1���wZ�o#D;��o6 ���U�Z�����۸I��Hﯲ��8�&{�)J/cME��Rg?��oO����(�t2�$R��7�2j�Y+���Ti��>	)�2��G��N]`��� �G*���U`j��x�F�?*͍��˹f��mlll����:�EdHn�������f'���Ni����4��|�M�}HG>���Z���TC����Vk��_{�$*Qx�k#�"��E��&G�e�ɒ��\����3�a]Ai��`����i���w��s�zy�~���XW�W2���,�lu�%�ᬨ�dLѓX�Z�����IG<�!�G����ٚ�/i1�7��Vd,��j�w�K@����B�5��U��ܽ������m��|,�Rk.v1[@�	�?����<�PK   �|�X��ί�  6'     jsons/user_defined.json�[o�6ǿ��3�/y����4+0%Q� Gre;AQ����'�DY̲�a����r��9��6\]���p�2���$if��hxg�U�g�`���&,_]����Ǚ�-��&���i�৙�#?�/"�6�y��~����[��ٺ�S?�*�d�>L�beF��^�D �@�B
#K�GI�#�ش�YEE�\��~��F��0F$��� 4
%P�D *.���@����~�|	K�n�+o�V�G�4�fI><�6�6��t�\�G����@��=>����3��W[��p��_6�q�4���Ԓ�`�/䫴��i�(�rIΰ�#DU�$G�l��q���|7d������]�s{:>9���b�}�NE]Tܓʮ�����=���%]о==�O���I��]�Ϗ/���۷���&^P�%P�3�.�h�Ò`�7a���xr0�;)�E�����ˏN�j"�?��Բ�PoF�zNF��A���9	-k���	>�O�nH�ڀ���̏Nܐ�� �C���Ӄ1ws��W�Vb܌����>�uW��Ի��t�o*�B�u7��T�Įj�r�M���}�`ͱˇ�T���'u�n
� ���AnP�����]�/qZ���k�Tq��в�s�.\M�܀������yܲ�S_@�^�[�u⋰���~˞}폙;~m�[y��n�MQ{�`L��r���|S����Ҕ�����*i����ǳ�wn@S�ޮO�:f�)_�������T�z?��4�O[�pY�KS��mb[�X��9w]��]fe�B/6Ui����3l��ú,p�ߟgG��r���q���pav�
�eS��V��vu�It���x�ޕ<�.�G�Y]�`F1ɱ��P%�*f@���EHe�:Fd9yf���C5YK��ڜ���I�r�9�э�������t6X�l��:�N���WW��"qj`84 3&��� �cˈ!\�Ƚ�7Q���C�FP#��� �J�(5����HCw��(�`��*������Q�RRu{�դ#�i��;먾b|_,2}�Qyu���m���_O���_�[L�xS~c���jE�r�B�"@m�B�B B"ca��2~S�Z����S�	V�l09����Ezg��|�^n�e+bi.`Bk ��QO��J`�����6��� b�]�C@!Mb�ed; ���HDB�0�%V�'	@ºf""�U�G�<PXAަ�'�|�OT@9�b�*�'=�p��ZJ��)���J���h�S���	����v0m,U��#�NO�	�(@S��|W�L��d�о�;r����QP�U$@�r���LK����]k%�ʑ{���"1��[�VցD�J�s v������>$i)j� �� ����@�S���Ĕ�0���}�_,�ѵb�$=!n嵜b�!�J�bJ�0�pyb�z��M��u�S�	FM ��Aj�b� ��-���D�.���[�-�xS����5#��lj�8�_DU�w�<�ׯI�BPt�__/�`~�����j�Z?���Y[@To�U<��B�����BAb��,�(I�	i�x(��FW�i}�FAF�4��U��L>�C��|H m���o#�/��m߰�fG�n'|D��m�dw�s����8�i��\����~ơ0PQ� a�*!2RvFQ���*J�t�o���Y��g}��PK
   �|�X�?p�Y  j�                   cirkitFile.jsonPK
   �l�XN|jo�  �  /             �  images/07e09445-3584-4801-8c96-91d92a49cf18.pngPK
   �|�X=A�'>    /             �   images/184639ba-f95c-4173-b99b-7b38d7e1948d.pngPK
   �|�X�wM�|  w  /             V<  images/5e95862a-04ad-4971-a9d5-8bbbb67b4e45.pngPK
   �|�X`$} [ /             X  images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK
   �|�X��O*�� ~� /             �� images/bd13d416-9901-4cb8-93ec-096849d17163.pngPK
   �|�X	� .W /             ��
 images/cca7adb9-3a17-4e0c-97e4-0d979b0e08a4.pngPK
   �|�X�+�s;  z;  /             ʿ images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK
   �l�X�4#�c  �  /             �� images/fa0dec76-8343-40ea-91a3-e67b9f04a458.pngPK
   �|�X��ί�  6'               �_ jsons/user_defined.jsonPK    
 
 j  yf   